library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity wallace_tree_24 is
    Port ( x : in STD_LOGIC_VECTOR (23 downto 0);
           y : in STD_LOGIC_VECTOR (23 downto 0);
           p : out STD_LOGIC_VECTOR (47 downto 0));
end wallace_tree_24;

architecture arch of wallace_tree_24 is

component carry_lookahead_adder_48 is
    Port ( x : in STD_LOGIC_VECTOR (47 downto 0);
           y : in STD_LOGIC_VECTOR (47 downto 0);
           cin : in STD_LOGIC;
           s : out STD_LOGIC_VECTOR (47 downto 0);
           cout : out STD_LOGIC);
end component;

component full_adder is
    Port ( x : in STD_LOGIC;
           y : in STD_LOGIC;
           cin : in STD_LOGIC;
           s : out STD_LOGIC;
           p : out STD_LOGIC;
           g : out STD_LOGIC;
           cout : out STD_LOGIC);
end component;

component half_adder is
    Port ( x : in STD_LOGIC;
           y : in STD_LOGIC;
           s : out STD_LOGIC;
           cout : out STD_LOGIC);
end component;

signal l1c0_0 : std_logic;
signal l1c1_0 : std_logic;
signal l1c1_1 : std_logic;
signal l1c2_0 : std_logic;
signal l1c2_1 : std_logic;
signal l1c2_2 : std_logic;
signal l1c3_0 : std_logic;
signal l1c3_1 : std_logic;
signal l1c3_2 : std_logic;
signal l1c3_3 : std_logic;
signal l1c4_0 : std_logic;
signal l1c4_1 : std_logic;
signal l1c4_2 : std_logic;
signal l1c4_3 : std_logic;
signal l1c4_4 : std_logic;
signal l1c5_0 : std_logic;
signal l1c5_1 : std_logic;
signal l1c5_2 : std_logic;
signal l1c5_3 : std_logic;
signal l1c5_4 : std_logic;
signal l1c5_5 : std_logic;
signal l1c6_0 : std_logic;
signal l1c6_1 : std_logic;
signal l1c6_2 : std_logic;
signal l1c6_3 : std_logic;
signal l1c6_4 : std_logic;
signal l1c6_5 : std_logic;
signal l1c6_6 : std_logic;
signal l1c7_0 : std_logic;
signal l1c7_1 : std_logic;
signal l1c7_2 : std_logic;
signal l1c7_3 : std_logic;
signal l1c7_4 : std_logic;
signal l1c7_5 : std_logic;
signal l1c7_6 : std_logic;
signal l1c7_7 : std_logic;
signal l1c8_0 : std_logic;
signal l1c8_1 : std_logic;
signal l1c8_2 : std_logic;
signal l1c8_3 : std_logic;
signal l1c8_4 : std_logic;
signal l1c8_5 : std_logic;
signal l1c8_6 : std_logic;
signal l1c8_7 : std_logic;
signal l1c8_8 : std_logic;
signal l1c9_0 : std_logic;
signal l1c9_1 : std_logic;
signal l1c9_2 : std_logic;
signal l1c9_3 : std_logic;
signal l1c9_4 : std_logic;
signal l1c9_5 : std_logic;
signal l1c9_6 : std_logic;
signal l1c9_7 : std_logic;
signal l1c9_8 : std_logic;
signal l1c9_9 : std_logic;
signal l1c10_0 : std_logic;
signal l1c10_1 : std_logic;
signal l1c10_2 : std_logic;
signal l1c10_3 : std_logic;
signal l1c10_4 : std_logic;
signal l1c10_5 : std_logic;
signal l1c10_6 : std_logic;
signal l1c10_7 : std_logic;
signal l1c10_8 : std_logic;
signal l1c10_9 : std_logic;
signal l1c10_10 : std_logic;
signal l1c11_0 : std_logic;
signal l1c11_1 : std_logic;
signal l1c11_2 : std_logic;
signal l1c11_3 : std_logic;
signal l1c11_4 : std_logic;
signal l1c11_5 : std_logic;
signal l1c11_6 : std_logic;
signal l1c11_7 : std_logic;
signal l1c11_8 : std_logic;
signal l1c11_9 : std_logic;
signal l1c11_10 : std_logic;
signal l1c11_11 : std_logic;
signal l1c12_0 : std_logic;
signal l1c12_1 : std_logic;
signal l1c12_2 : std_logic;
signal l1c12_3 : std_logic;
signal l1c12_4 : std_logic;
signal l1c12_5 : std_logic;
signal l1c12_6 : std_logic;
signal l1c12_7 : std_logic;
signal l1c12_8 : std_logic;
signal l1c12_9 : std_logic;
signal l1c12_10 : std_logic;
signal l1c12_11 : std_logic;
signal l1c12_12 : std_logic;
signal l1c13_0 : std_logic;
signal l1c13_1 : std_logic;
signal l1c13_2 : std_logic;
signal l1c13_3 : std_logic;
signal l1c13_4 : std_logic;
signal l1c13_5 : std_logic;
signal l1c13_6 : std_logic;
signal l1c13_7 : std_logic;
signal l1c13_8 : std_logic;
signal l1c13_9 : std_logic;
signal l1c13_10 : std_logic;
signal l1c13_11 : std_logic;
signal l1c13_12 : std_logic;
signal l1c13_13 : std_logic;
signal l1c14_0 : std_logic;
signal l1c14_1 : std_logic;
signal l1c14_2 : std_logic;
signal l1c14_3 : std_logic;
signal l1c14_4 : std_logic;
signal l1c14_5 : std_logic;
signal l1c14_6 : std_logic;
signal l1c14_7 : std_logic;
signal l1c14_8 : std_logic;
signal l1c14_9 : std_logic;
signal l1c14_10 : std_logic;
signal l1c14_11 : std_logic;
signal l1c14_12 : std_logic;
signal l1c14_13 : std_logic;
signal l1c14_14 : std_logic;
signal l1c15_0 : std_logic;
signal l1c15_1 : std_logic;
signal l1c15_2 : std_logic;
signal l1c15_3 : std_logic;
signal l1c15_4 : std_logic;
signal l1c15_5 : std_logic;
signal l1c15_6 : std_logic;
signal l1c15_7 : std_logic;
signal l1c15_8 : std_logic;
signal l1c15_9 : std_logic;
signal l1c15_10 : std_logic;
signal l1c15_11 : std_logic;
signal l1c15_12 : std_logic;
signal l1c15_13 : std_logic;
signal l1c15_14 : std_logic;
signal l1c15_15 : std_logic;
signal l1c16_0 : std_logic;
signal l1c16_1 : std_logic;
signal l1c16_2 : std_logic;
signal l1c16_3 : std_logic;
signal l1c16_4 : std_logic;
signal l1c16_5 : std_logic;
signal l1c16_6 : std_logic;
signal l1c16_7 : std_logic;
signal l1c16_8 : std_logic;
signal l1c16_9 : std_logic;
signal l1c16_10 : std_logic;
signal l1c16_11 : std_logic;
signal l1c16_12 : std_logic;
signal l1c16_13 : std_logic;
signal l1c16_14 : std_logic;
signal l1c16_15 : std_logic;
signal l1c16_16 : std_logic;
signal l1c17_0 : std_logic;
signal l1c17_1 : std_logic;
signal l1c17_2 : std_logic;
signal l1c17_3 : std_logic;
signal l1c17_4 : std_logic;
signal l1c17_5 : std_logic;
signal l1c17_6 : std_logic;
signal l1c17_7 : std_logic;
signal l1c17_8 : std_logic;
signal l1c17_9 : std_logic;
signal l1c17_10 : std_logic;
signal l1c17_11 : std_logic;
signal l1c17_12 : std_logic;
signal l1c17_13 : std_logic;
signal l1c17_14 : std_logic;
signal l1c17_15 : std_logic;
signal l1c17_16 : std_logic;
signal l1c17_17 : std_logic;
signal l1c18_0 : std_logic;
signal l1c18_1 : std_logic;
signal l1c18_2 : std_logic;
signal l1c18_3 : std_logic;
signal l1c18_4 : std_logic;
signal l1c18_5 : std_logic;
signal l1c18_6 : std_logic;
signal l1c18_7 : std_logic;
signal l1c18_8 : std_logic;
signal l1c18_9 : std_logic;
signal l1c18_10 : std_logic;
signal l1c18_11 : std_logic;
signal l1c18_12 : std_logic;
signal l1c18_13 : std_logic;
signal l1c18_14 : std_logic;
signal l1c18_15 : std_logic;
signal l1c18_16 : std_logic;
signal l1c18_17 : std_logic;
signal l1c18_18 : std_logic;
signal l1c19_0 : std_logic;
signal l1c19_1 : std_logic;
signal l1c19_2 : std_logic;
signal l1c19_3 : std_logic;
signal l1c19_4 : std_logic;
signal l1c19_5 : std_logic;
signal l1c19_6 : std_logic;
signal l1c19_7 : std_logic;
signal l1c19_8 : std_logic;
signal l1c19_9 : std_logic;
signal l1c19_10 : std_logic;
signal l1c19_11 : std_logic;
signal l1c19_12 : std_logic;
signal l1c19_13 : std_logic;
signal l1c19_14 : std_logic;
signal l1c19_15 : std_logic;
signal l1c19_16 : std_logic;
signal l1c19_17 : std_logic;
signal l1c19_18 : std_logic;
signal l1c19_19 : std_logic;
signal l1c20_0 : std_logic;
signal l1c20_1 : std_logic;
signal l1c20_2 : std_logic;
signal l1c20_3 : std_logic;
signal l1c20_4 : std_logic;
signal l1c20_5 : std_logic;
signal l1c20_6 : std_logic;
signal l1c20_7 : std_logic;
signal l1c20_8 : std_logic;
signal l1c20_9 : std_logic;
signal l1c20_10 : std_logic;
signal l1c20_11 : std_logic;
signal l1c20_12 : std_logic;
signal l1c20_13 : std_logic;
signal l1c20_14 : std_logic;
signal l1c20_15 : std_logic;
signal l1c20_16 : std_logic;
signal l1c20_17 : std_logic;
signal l1c20_18 : std_logic;
signal l1c20_19 : std_logic;
signal l1c20_20 : std_logic;
signal l1c21_0 : std_logic;
signal l1c21_1 : std_logic;
signal l1c21_2 : std_logic;
signal l1c21_3 : std_logic;
signal l1c21_4 : std_logic;
signal l1c21_5 : std_logic;
signal l1c21_6 : std_logic;
signal l1c21_7 : std_logic;
signal l1c21_8 : std_logic;
signal l1c21_9 : std_logic;
signal l1c21_10 : std_logic;
signal l1c21_11 : std_logic;
signal l1c21_12 : std_logic;
signal l1c21_13 : std_logic;
signal l1c21_14 : std_logic;
signal l1c21_15 : std_logic;
signal l1c21_16 : std_logic;
signal l1c21_17 : std_logic;
signal l1c21_18 : std_logic;
signal l1c21_19 : std_logic;
signal l1c21_20 : std_logic;
signal l1c21_21 : std_logic;
signal l1c22_0 : std_logic;
signal l1c22_1 : std_logic;
signal l1c22_2 : std_logic;
signal l1c22_3 : std_logic;
signal l1c22_4 : std_logic;
signal l1c22_5 : std_logic;
signal l1c22_6 : std_logic;
signal l1c22_7 : std_logic;
signal l1c22_8 : std_logic;
signal l1c22_9 : std_logic;
signal l1c22_10 : std_logic;
signal l1c22_11 : std_logic;
signal l1c22_12 : std_logic;
signal l1c22_13 : std_logic;
signal l1c22_14 : std_logic;
signal l1c22_15 : std_logic;
signal l1c22_16 : std_logic;
signal l1c22_17 : std_logic;
signal l1c22_18 : std_logic;
signal l1c22_19 : std_logic;
signal l1c22_20 : std_logic;
signal l1c22_21 : std_logic;
signal l1c22_22 : std_logic;
signal l1c23_0 : std_logic;
signal l1c23_1 : std_logic;
signal l1c23_2 : std_logic;
signal l1c23_3 : std_logic;
signal l1c23_4 : std_logic;
signal l1c23_5 : std_logic;
signal l1c23_6 : std_logic;
signal l1c23_7 : std_logic;
signal l1c23_8 : std_logic;
signal l1c23_9 : std_logic;
signal l1c23_10 : std_logic;
signal l1c23_11 : std_logic;
signal l1c23_12 : std_logic;
signal l1c23_13 : std_logic;
signal l1c23_14 : std_logic;
signal l1c23_15 : std_logic;
signal l1c23_16 : std_logic;
signal l1c23_17 : std_logic;
signal l1c23_18 : std_logic;
signal l1c23_19 : std_logic;
signal l1c23_20 : std_logic;
signal l1c23_21 : std_logic;
signal l1c23_22 : std_logic;
signal l1c23_23 : std_logic;
signal l1c24_0 : std_logic;
signal l1c24_1 : std_logic;
signal l1c24_2 : std_logic;
signal l1c24_3 : std_logic;
signal l1c24_4 : std_logic;
signal l1c24_5 : std_logic;
signal l1c24_6 : std_logic;
signal l1c24_7 : std_logic;
signal l1c24_8 : std_logic;
signal l1c24_9 : std_logic;
signal l1c24_10 : std_logic;
signal l1c24_11 : std_logic;
signal l1c24_12 : std_logic;
signal l1c24_13 : std_logic;
signal l1c24_14 : std_logic;
signal l1c24_15 : std_logic;
signal l1c24_16 : std_logic;
signal l1c24_17 : std_logic;
signal l1c24_18 : std_logic;
signal l1c24_19 : std_logic;
signal l1c24_20 : std_logic;
signal l1c24_21 : std_logic;
signal l1c24_22 : std_logic;
signal l1c25_0 : std_logic;
signal l1c25_1 : std_logic;
signal l1c25_2 : std_logic;
signal l1c25_3 : std_logic;
signal l1c25_4 : std_logic;
signal l1c25_5 : std_logic;
signal l1c25_6 : std_logic;
signal l1c25_7 : std_logic;
signal l1c25_8 : std_logic;
signal l1c25_9 : std_logic;
signal l1c25_10 : std_logic;
signal l1c25_11 : std_logic;
signal l1c25_12 : std_logic;
signal l1c25_13 : std_logic;
signal l1c25_14 : std_logic;
signal l1c25_15 : std_logic;
signal l1c25_16 : std_logic;
signal l1c25_17 : std_logic;
signal l1c25_18 : std_logic;
signal l1c25_19 : std_logic;
signal l1c25_20 : std_logic;
signal l1c25_21 : std_logic;
signal l1c26_0 : std_logic;
signal l1c26_1 : std_logic;
signal l1c26_2 : std_logic;
signal l1c26_3 : std_logic;
signal l1c26_4 : std_logic;
signal l1c26_5 : std_logic;
signal l1c26_6 : std_logic;
signal l1c26_7 : std_logic;
signal l1c26_8 : std_logic;
signal l1c26_9 : std_logic;
signal l1c26_10 : std_logic;
signal l1c26_11 : std_logic;
signal l1c26_12 : std_logic;
signal l1c26_13 : std_logic;
signal l1c26_14 : std_logic;
signal l1c26_15 : std_logic;
signal l1c26_16 : std_logic;
signal l1c26_17 : std_logic;
signal l1c26_18 : std_logic;
signal l1c26_19 : std_logic;
signal l1c26_20 : std_logic;
signal l1c27_0 : std_logic;
signal l1c27_1 : std_logic;
signal l1c27_2 : std_logic;
signal l1c27_3 : std_logic;
signal l1c27_4 : std_logic;
signal l1c27_5 : std_logic;
signal l1c27_6 : std_logic;
signal l1c27_7 : std_logic;
signal l1c27_8 : std_logic;
signal l1c27_9 : std_logic;
signal l1c27_10 : std_logic;
signal l1c27_11 : std_logic;
signal l1c27_12 : std_logic;
signal l1c27_13 : std_logic;
signal l1c27_14 : std_logic;
signal l1c27_15 : std_logic;
signal l1c27_16 : std_logic;
signal l1c27_17 : std_logic;
signal l1c27_18 : std_logic;
signal l1c27_19 : std_logic;
signal l1c28_0 : std_logic;
signal l1c28_1 : std_logic;
signal l1c28_2 : std_logic;
signal l1c28_3 : std_logic;
signal l1c28_4 : std_logic;
signal l1c28_5 : std_logic;
signal l1c28_6 : std_logic;
signal l1c28_7 : std_logic;
signal l1c28_8 : std_logic;
signal l1c28_9 : std_logic;
signal l1c28_10 : std_logic;
signal l1c28_11 : std_logic;
signal l1c28_12 : std_logic;
signal l1c28_13 : std_logic;
signal l1c28_14 : std_logic;
signal l1c28_15 : std_logic;
signal l1c28_16 : std_logic;
signal l1c28_17 : std_logic;
signal l1c28_18 : std_logic;
signal l1c29_0 : std_logic;
signal l1c29_1 : std_logic;
signal l1c29_2 : std_logic;
signal l1c29_3 : std_logic;
signal l1c29_4 : std_logic;
signal l1c29_5 : std_logic;
signal l1c29_6 : std_logic;
signal l1c29_7 : std_logic;
signal l1c29_8 : std_logic;
signal l1c29_9 : std_logic;
signal l1c29_10 : std_logic;
signal l1c29_11 : std_logic;
signal l1c29_12 : std_logic;
signal l1c29_13 : std_logic;
signal l1c29_14 : std_logic;
signal l1c29_15 : std_logic;
signal l1c29_16 : std_logic;
signal l1c29_17 : std_logic;
signal l1c30_0 : std_logic;
signal l1c30_1 : std_logic;
signal l1c30_2 : std_logic;
signal l1c30_3 : std_logic;
signal l1c30_4 : std_logic;
signal l1c30_5 : std_logic;
signal l1c30_6 : std_logic;
signal l1c30_7 : std_logic;
signal l1c30_8 : std_logic;
signal l1c30_9 : std_logic;
signal l1c30_10 : std_logic;
signal l1c30_11 : std_logic;
signal l1c30_12 : std_logic;
signal l1c30_13 : std_logic;
signal l1c30_14 : std_logic;
signal l1c30_15 : std_logic;
signal l1c30_16 : std_logic;
signal l1c31_0 : std_logic;
signal l1c31_1 : std_logic;
signal l1c31_2 : std_logic;
signal l1c31_3 : std_logic;
signal l1c31_4 : std_logic;
signal l1c31_5 : std_logic;
signal l1c31_6 : std_logic;
signal l1c31_7 : std_logic;
signal l1c31_8 : std_logic;
signal l1c31_9 : std_logic;
signal l1c31_10 : std_logic;
signal l1c31_11 : std_logic;
signal l1c31_12 : std_logic;
signal l1c31_13 : std_logic;
signal l1c31_14 : std_logic;
signal l1c31_15 : std_logic;
signal l1c32_0 : std_logic;
signal l1c32_1 : std_logic;
signal l1c32_2 : std_logic;
signal l1c32_3 : std_logic;
signal l1c32_4 : std_logic;
signal l1c32_5 : std_logic;
signal l1c32_6 : std_logic;
signal l1c32_7 : std_logic;
signal l1c32_8 : std_logic;
signal l1c32_9 : std_logic;
signal l1c32_10 : std_logic;
signal l1c32_11 : std_logic;
signal l1c32_12 : std_logic;
signal l1c32_13 : std_logic;
signal l1c32_14 : std_logic;
signal l1c33_0 : std_logic;
signal l1c33_1 : std_logic;
signal l1c33_2 : std_logic;
signal l1c33_3 : std_logic;
signal l1c33_4 : std_logic;
signal l1c33_5 : std_logic;
signal l1c33_6 : std_logic;
signal l1c33_7 : std_logic;
signal l1c33_8 : std_logic;
signal l1c33_9 : std_logic;
signal l1c33_10 : std_logic;
signal l1c33_11 : std_logic;
signal l1c33_12 : std_logic;
signal l1c33_13 : std_logic;
signal l1c34_0 : std_logic;
signal l1c34_1 : std_logic;
signal l1c34_2 : std_logic;
signal l1c34_3 : std_logic;
signal l1c34_4 : std_logic;
signal l1c34_5 : std_logic;
signal l1c34_6 : std_logic;
signal l1c34_7 : std_logic;
signal l1c34_8 : std_logic;
signal l1c34_9 : std_logic;
signal l1c34_10 : std_logic;
signal l1c34_11 : std_logic;
signal l1c34_12 : std_logic;
signal l1c35_0 : std_logic;
signal l1c35_1 : std_logic;
signal l1c35_2 : std_logic;
signal l1c35_3 : std_logic;
signal l1c35_4 : std_logic;
signal l1c35_5 : std_logic;
signal l1c35_6 : std_logic;
signal l1c35_7 : std_logic;
signal l1c35_8 : std_logic;
signal l1c35_9 : std_logic;
signal l1c35_10 : std_logic;
signal l1c35_11 : std_logic;
signal l1c36_0 : std_logic;
signal l1c36_1 : std_logic;
signal l1c36_2 : std_logic;
signal l1c36_3 : std_logic;
signal l1c36_4 : std_logic;
signal l1c36_5 : std_logic;
signal l1c36_6 : std_logic;
signal l1c36_7 : std_logic;
signal l1c36_8 : std_logic;
signal l1c36_9 : std_logic;
signal l1c36_10 : std_logic;
signal l1c37_0 : std_logic;
signal l1c37_1 : std_logic;
signal l1c37_2 : std_logic;
signal l1c37_3 : std_logic;
signal l1c37_4 : std_logic;
signal l1c37_5 : std_logic;
signal l1c37_6 : std_logic;
signal l1c37_7 : std_logic;
signal l1c37_8 : std_logic;
signal l1c37_9 : std_logic;
signal l1c38_0 : std_logic;
signal l1c38_1 : std_logic;
signal l1c38_2 : std_logic;
signal l1c38_3 : std_logic;
signal l1c38_4 : std_logic;
signal l1c38_5 : std_logic;
signal l1c38_6 : std_logic;
signal l1c38_7 : std_logic;
signal l1c38_8 : std_logic;
signal l1c39_0 : std_logic;
signal l1c39_1 : std_logic;
signal l1c39_2 : std_logic;
signal l1c39_3 : std_logic;
signal l1c39_4 : std_logic;
signal l1c39_5 : std_logic;
signal l1c39_6 : std_logic;
signal l1c39_7 : std_logic;
signal l1c40_0 : std_logic;
signal l1c40_1 : std_logic;
signal l1c40_2 : std_logic;
signal l1c40_3 : std_logic;
signal l1c40_4 : std_logic;
signal l1c40_5 : std_logic;
signal l1c40_6 : std_logic;
signal l1c41_0 : std_logic;
signal l1c41_1 : std_logic;
signal l1c41_2 : std_logic;
signal l1c41_3 : std_logic;
signal l1c41_4 : std_logic;
signal l1c41_5 : std_logic;
signal l1c42_0 : std_logic;
signal l1c42_1 : std_logic;
signal l1c42_2 : std_logic;
signal l1c42_3 : std_logic;
signal l1c42_4 : std_logic;
signal l1c43_0 : std_logic;
signal l1c43_1 : std_logic;
signal l1c43_2 : std_logic;
signal l1c43_3 : std_logic;
signal l1c44_0 : std_logic;
signal l1c44_1 : std_logic;
signal l1c44_2 : std_logic;
signal l1c45_0 : std_logic;
signal l1c45_1 : std_logic;
signal l1c46_0 : std_logic;
signal l2c1_0 : std_logic;
signal l2c2_0 : std_logic;
signal l2c2_1 : std_logic;
signal l2c3_0 : std_logic;
signal l2c3_1 : std_logic;
signal l2c4_0 : std_logic;
signal l2c4_1 : std_logic;
signal l2c5_0 : std_logic;
signal l2c4_2 : std_logic;
signal l2c5_1 : std_logic;
signal l2c5_2 : std_logic;
signal l2c6_0 : std_logic;
signal l2c5_3 : std_logic;
signal l2c6_1 : std_logic;
signal l2c6_2 : std_logic;
signal l2c7_0 : std_logic;
signal l2c6_3 : std_logic;
signal l2c7_1 : std_logic;
signal l2c7_2 : std_logic;
signal l2c8_0 : std_logic;
signal l2c7_3 : std_logic;
signal l2c8_1 : std_logic;
signal l2c7_4 : std_logic;
signal l2c8_2 : std_logic;
signal l2c8_3 : std_logic;
signal l2c9_0 : std_logic;
signal l2c8_4 : std_logic;
signal l2c9_1 : std_logic;
signal l2c8_5 : std_logic;
signal l2c9_2 : std_logic;
signal l2c9_3 : std_logic;
signal l2c10_0 : std_logic;
signal l2c9_4 : std_logic;
signal l2c10_1 : std_logic;
signal l2c9_5 : std_logic;
signal l2c10_2 : std_logic;
signal l2c10_3 : std_logic;
signal l2c11_0 : std_logic;
signal l2c10_4 : std_logic;
signal l2c11_1 : std_logic;
signal l2c10_5 : std_logic;
signal l2c11_2 : std_logic;
signal l2c10_6 : std_logic;
signal l2c11_3 : std_logic;
signal l2c11_4 : std_logic;
signal l2c12_0 : std_logic;
signal l2c11_5 : std_logic;
signal l2c12_1 : std_logic;
signal l2c11_6 : std_logic;
signal l2c12_2 : std_logic;
signal l2c11_7 : std_logic;
signal l2c12_3 : std_logic;
signal l2c12_4 : std_logic;
signal l2c13_0 : std_logic;
signal l2c12_5 : std_logic;
signal l2c13_1 : std_logic;
signal l2c12_6 : std_logic;
signal l2c13_2 : std_logic;
signal l2c12_7 : std_logic;
signal l2c13_3 : std_logic;
signal l2c13_4 : std_logic;
signal l2c14_0 : std_logic;
signal l2c13_5 : std_logic;
signal l2c14_1 : std_logic;
signal l2c13_6 : std_logic;
signal l2c14_2 : std_logic;
signal l2c13_7 : std_logic;
signal l2c14_3 : std_logic;
signal l2c13_8 : std_logic;
signal l2c14_4 : std_logic;
signal l2c14_5 : std_logic;
signal l2c15_0 : std_logic;
signal l2c14_6 : std_logic;
signal l2c15_1 : std_logic;
signal l2c14_7 : std_logic;
signal l2c15_2 : std_logic;
signal l2c14_8 : std_logic;
signal l2c15_3 : std_logic;
signal l2c14_9 : std_logic;
signal l2c15_4 : std_logic;
signal l2c15_5 : std_logic;
signal l2c16_0 : std_logic;
signal l2c15_6 : std_logic;
signal l2c16_1 : std_logic;
signal l2c15_7 : std_logic;
signal l2c16_2 : std_logic;
signal l2c15_8 : std_logic;
signal l2c16_3 : std_logic;
signal l2c15_9 : std_logic;
signal l2c16_4 : std_logic;
signal l2c16_5 : std_logic;
signal l2c17_0 : std_logic;
signal l2c16_6 : std_logic;
signal l2c17_1 : std_logic;
signal l2c16_7 : std_logic;
signal l2c17_2 : std_logic;
signal l2c16_8 : std_logic;
signal l2c17_3 : std_logic;
signal l2c16_9 : std_logic;
signal l2c17_4 : std_logic;
signal l2c16_10 : std_logic;
signal l2c17_5 : std_logic;
signal l2c17_6 : std_logic;
signal l2c18_0 : std_logic;
signal l2c17_7 : std_logic;
signal l2c18_1 : std_logic;
signal l2c17_8 : std_logic;
signal l2c18_2 : std_logic;
signal l2c17_9 : std_logic;
signal l2c18_3 : std_logic;
signal l2c17_10 : std_logic;
signal l2c18_4 : std_logic;
signal l2c17_11 : std_logic;
signal l2c18_5 : std_logic;
signal l2c18_6 : std_logic;
signal l2c19_0 : std_logic;
signal l2c18_7 : std_logic;
signal l2c19_1 : std_logic;
signal l2c18_8 : std_logic;
signal l2c19_2 : std_logic;
signal l2c18_9 : std_logic;
signal l2c19_3 : std_logic;
signal l2c18_10 : std_logic;
signal l2c19_4 : std_logic;
signal l2c18_11 : std_logic;
signal l2c19_5 : std_logic;
signal l2c19_6 : std_logic;
signal l2c20_0 : std_logic;
signal l2c19_7 : std_logic;
signal l2c20_1 : std_logic;
signal l2c19_8 : std_logic;
signal l2c20_2 : std_logic;
signal l2c19_9 : std_logic;
signal l2c20_3 : std_logic;
signal l2c19_10 : std_logic;
signal l2c20_4 : std_logic;
signal l2c19_11 : std_logic;
signal l2c20_5 : std_logic;
signal l2c19_12 : std_logic;
signal l2c20_6 : std_logic;
signal l2c20_7 : std_logic;
signal l2c21_0 : std_logic;
signal l2c20_8 : std_logic;
signal l2c21_1 : std_logic;
signal l2c20_9 : std_logic;
signal l2c21_2 : std_logic;
signal l2c20_10 : std_logic;
signal l2c21_3 : std_logic;
signal l2c20_11 : std_logic;
signal l2c21_4 : std_logic;
signal l2c20_12 : std_logic;
signal l2c21_5 : std_logic;
signal l2c20_13 : std_logic;
signal l2c21_6 : std_logic;
signal l2c21_7 : std_logic;
signal l2c22_0 : std_logic;
signal l2c21_8 : std_logic;
signal l2c22_1 : std_logic;
signal l2c21_9 : std_logic;
signal l2c22_2 : std_logic;
signal l2c21_10 : std_logic;
signal l2c22_3 : std_logic;
signal l2c21_11 : std_logic;
signal l2c22_4 : std_logic;
signal l2c21_12 : std_logic;
signal l2c22_5 : std_logic;
signal l2c21_13 : std_logic;
signal l2c22_6 : std_logic;
signal l2c22_7 : std_logic;
signal l2c23_0 : std_logic;
signal l2c22_8 : std_logic;
signal l2c23_1 : std_logic;
signal l2c22_9 : std_logic;
signal l2c23_2 : std_logic;
signal l2c22_10 : std_logic;
signal l2c23_3 : std_logic;
signal l2c22_11 : std_logic;
signal l2c23_4 : std_logic;
signal l2c22_12 : std_logic;
signal l2c23_5 : std_logic;
signal l2c22_13 : std_logic;
signal l2c23_6 : std_logic;
signal l2c22_14 : std_logic;
signal l2c23_7 : std_logic;
signal l2c23_8 : std_logic;
signal l2c24_0 : std_logic;
signal l2c23_9 : std_logic;
signal l2c24_1 : std_logic;
signal l2c23_10 : std_logic;
signal l2c24_2 : std_logic;
signal l2c23_11 : std_logic;
signal l2c24_3 : std_logic;
signal l2c23_12 : std_logic;
signal l2c24_4 : std_logic;
signal l2c23_13 : std_logic;
signal l2c24_5 : std_logic;
signal l2c23_14 : std_logic;
signal l2c24_6 : std_logic;
signal l2c23_15 : std_logic;
signal l2c24_7 : std_logic;
signal l2c24_8 : std_logic;
signal l2c25_0 : std_logic;
signal l2c24_9 : std_logic;
signal l2c25_1 : std_logic;
signal l2c24_10 : std_logic;
signal l2c25_2 : std_logic;
signal l2c24_11 : std_logic;
signal l2c25_3 : std_logic;
signal l2c24_12 : std_logic;
signal l2c25_4 : std_logic;
signal l2c24_13 : std_logic;
signal l2c25_5 : std_logic;
signal l2c24_14 : std_logic;
signal l2c25_6 : std_logic;
signal l2c24_15 : std_logic;
signal l2c25_7 : std_logic;
signal l2c25_8 : std_logic;
signal l2c26_0 : std_logic;
signal l2c25_9 : std_logic;
signal l2c26_1 : std_logic;
signal l2c25_10 : std_logic;
signal l2c26_2 : std_logic;
signal l2c25_11 : std_logic;
signal l2c26_3 : std_logic;
signal l2c25_12 : std_logic;
signal l2c26_4 : std_logic;
signal l2c25_13 : std_logic;
signal l2c26_5 : std_logic;
signal l2c25_14 : std_logic;
signal l2c26_6 : std_logic;
signal l2c26_7 : std_logic;
signal l2c27_0 : std_logic;
signal l2c26_8 : std_logic;
signal l2c27_1 : std_logic;
signal l2c26_9 : std_logic;
signal l2c27_2 : std_logic;
signal l2c26_10 : std_logic;
signal l2c27_3 : std_logic;
signal l2c26_11 : std_logic;
signal l2c27_4 : std_logic;
signal l2c26_12 : std_logic;
signal l2c27_5 : std_logic;
signal l2c26_13 : std_logic;
signal l2c27_6 : std_logic;
signal l2c27_7 : std_logic;
signal l2c28_0 : std_logic;
signal l2c27_8 : std_logic;
signal l2c28_1 : std_logic;
signal l2c27_9 : std_logic;
signal l2c28_2 : std_logic;
signal l2c27_10 : std_logic;
signal l2c28_3 : std_logic;
signal l2c27_11 : std_logic;
signal l2c28_4 : std_logic;
signal l2c27_12 : std_logic;
signal l2c28_5 : std_logic;
signal l2c27_13 : std_logic;
signal l2c28_6 : std_logic;
signal l2c28_7 : std_logic;
signal l2c29_0 : std_logic;
signal l2c28_8 : std_logic;
signal l2c29_1 : std_logic;
signal l2c28_9 : std_logic;
signal l2c29_2 : std_logic;
signal l2c28_10 : std_logic;
signal l2c29_3 : std_logic;
signal l2c28_11 : std_logic;
signal l2c29_4 : std_logic;
signal l2c28_12 : std_logic;
signal l2c29_5 : std_logic;
signal l2c29_6 : std_logic;
signal l2c30_0 : std_logic;
signal l2c29_7 : std_logic;
signal l2c30_1 : std_logic;
signal l2c29_8 : std_logic;
signal l2c30_2 : std_logic;
signal l2c29_9 : std_logic;
signal l2c30_3 : std_logic;
signal l2c29_10 : std_logic;
signal l2c30_4 : std_logic;
signal l2c29_11 : std_logic;
signal l2c30_5 : std_logic;
signal l2c30_6 : std_logic;
signal l2c31_0 : std_logic;
signal l2c30_7 : std_logic;
signal l2c31_1 : std_logic;
signal l2c30_8 : std_logic;
signal l2c31_2 : std_logic;
signal l2c30_9 : std_logic;
signal l2c31_3 : std_logic;
signal l2c30_10 : std_logic;
signal l2c31_4 : std_logic;
signal l2c30_11 : std_logic;
signal l2c31_5 : std_logic;
signal l2c31_6 : std_logic;
signal l2c32_0 : std_logic;
signal l2c31_7 : std_logic;
signal l2c32_1 : std_logic;
signal l2c31_8 : std_logic;
signal l2c32_2 : std_logic;
signal l2c31_9 : std_logic;
signal l2c32_3 : std_logic;
signal l2c31_10 : std_logic;
signal l2c32_4 : std_logic;
signal l2c32_5 : std_logic;
signal l2c33_0 : std_logic;
signal l2c32_6 : std_logic;
signal l2c33_1 : std_logic;
signal l2c32_7 : std_logic;
signal l2c33_2 : std_logic;
signal l2c32_8 : std_logic;
signal l2c33_3 : std_logic;
signal l2c32_9 : std_logic;
signal l2c33_4 : std_logic;
signal l2c33_5 : std_logic;
signal l2c34_0 : std_logic;
signal l2c33_6 : std_logic;
signal l2c34_1 : std_logic;
signal l2c33_7 : std_logic;
signal l2c34_2 : std_logic;
signal l2c33_8 : std_logic;
signal l2c34_3 : std_logic;
signal l2c33_9 : std_logic;
signal l2c34_4 : std_logic;
signal l2c34_5 : std_logic;
signal l2c35_0 : std_logic;
signal l2c34_6 : std_logic;
signal l2c35_1 : std_logic;
signal l2c34_7 : std_logic;
signal l2c35_2 : std_logic;
signal l2c34_8 : std_logic;
signal l2c35_3 : std_logic;
signal l2c35_4 : std_logic;
signal l2c36_0 : std_logic;
signal l2c35_5 : std_logic;
signal l2c36_1 : std_logic;
signal l2c35_6 : std_logic;
signal l2c36_2 : std_logic;
signal l2c35_7 : std_logic;
signal l2c36_3 : std_logic;
signal l2c36_4 : std_logic;
signal l2c37_0 : std_logic;
signal l2c36_5 : std_logic;
signal l2c37_1 : std_logic;
signal l2c36_6 : std_logic;
signal l2c37_2 : std_logic;
signal l2c36_7 : std_logic;
signal l2c37_3 : std_logic;
signal l2c37_4 : std_logic;
signal l2c38_0 : std_logic;
signal l2c37_5 : std_logic;
signal l2c38_1 : std_logic;
signal l2c37_6 : std_logic;
signal l2c38_2 : std_logic;
signal l2c38_3 : std_logic;
signal l2c39_0 : std_logic;
signal l2c38_4 : std_logic;
signal l2c39_1 : std_logic;
signal l2c38_5 : std_logic;
signal l2c39_2 : std_logic;
signal l2c39_3 : std_logic;
signal l2c40_0 : std_logic;
signal l2c39_4 : std_logic;
signal l2c40_1 : std_logic;
signal l2c39_5 : std_logic;
signal l2c40_2 : std_logic;
signal l2c40_3 : std_logic;
signal l2c41_0 : std_logic;
signal l2c40_4 : std_logic;
signal l2c41_1 : std_logic;
signal l2c41_2 : std_logic;
signal l2c42_0 : std_logic;
signal l2c41_3 : std_logic;
signal l2c42_1 : std_logic;
signal l2c42_2 : std_logic;
signal l2c43_0 : std_logic;
signal l2c42_3 : std_logic;
signal l2c43_1 : std_logic;
signal l2c43_2 : std_logic;
signal l2c44_0 : std_logic;
signal l2c44_1 : std_logic;
signal l2c45_0 : std_logic;
signal l2c45_1 : std_logic;
signal l2c46_0 : std_logic;
signal l3c2_0 : std_logic;
signal l3c3_0 : std_logic;
signal l3c3_1 : std_logic;
signal l3c4_0 : std_logic;
signal l3c4_1 : std_logic;
signal l3c5_0 : std_logic;
signal l3c5_1 : std_logic;
signal l3c6_0 : std_logic;
signal l3c6_1 : std_logic;
signal l3c7_0 : std_logic;
signal l3c6_2 : std_logic;
signal l3c7_1 : std_logic;
signal l3c7_2 : std_logic;
signal l3c8_0 : std_logic;
signal l3c7_3 : std_logic;
signal l3c8_1 : std_logic;
signal l3c8_2 : std_logic;
signal l3c9_0 : std_logic;
signal l3c8_3 : std_logic;
signal l3c9_1 : std_logic;
signal l3c9_2 : std_logic;
signal l3c10_0 : std_logic;
signal l3c9_3 : std_logic;
signal l3c10_1 : std_logic;
signal l3c10_2 : std_logic;
signal l3c11_0 : std_logic;
signal l3c10_3 : std_logic;
signal l3c11_1 : std_logic;
signal l3c11_2 : std_logic;
signal l3c12_0 : std_logic;
signal l3c11_3 : std_logic;
signal l3c12_1 : std_logic;
signal l3c11_4 : std_logic;
signal l3c12_2 : std_logic;
signal l3c12_3 : std_logic;
signal l3c13_0 : std_logic;
signal l3c12_4 : std_logic;
signal l3c13_1 : std_logic;
signal l3c12_5 : std_logic;
signal l3c13_2 : std_logic;
signal l3c13_3 : std_logic;
signal l3c14_0 : std_logic;
signal l3c13_4 : std_logic;
signal l3c14_1 : std_logic;
signal l3c13_5 : std_logic;
signal l3c14_2 : std_logic;
signal l3c14_3 : std_logic;
signal l3c15_0 : std_logic;
signal l3c14_4 : std_logic;
signal l3c15_1 : std_logic;
signal l3c14_5 : std_logic;
signal l3c15_2 : std_logic;
signal l3c15_3 : std_logic;
signal l3c16_0 : std_logic;
signal l3c15_4 : std_logic;
signal l3c16_1 : std_logic;
signal l3c15_5 : std_logic;
signal l3c16_2 : std_logic;
signal l3c15_6 : std_logic;
signal l3c16_3 : std_logic;
signal l3c16_4 : std_logic;
signal l3c17_0 : std_logic;
signal l3c16_5 : std_logic;
signal l3c17_1 : std_logic;
signal l3c16_6 : std_logic;
signal l3c17_2 : std_logic;
signal l3c16_7 : std_logic;
signal l3c17_3 : std_logic;
signal l3c17_4 : std_logic;
signal l3c18_0 : std_logic;
signal l3c17_5 : std_logic;
signal l3c18_1 : std_logic;
signal l3c17_6 : std_logic;
signal l3c18_2 : std_logic;
signal l3c17_7 : std_logic;
signal l3c18_3 : std_logic;
signal l3c18_4 : std_logic;
signal l3c19_0 : std_logic;
signal l3c18_5 : std_logic;
signal l3c19_1 : std_logic;
signal l3c18_6 : std_logic;
signal l3c19_2 : std_logic;
signal l3c18_7 : std_logic;
signal l3c19_3 : std_logic;
signal l3c19_4 : std_logic;
signal l3c20_0 : std_logic;
signal l3c19_5 : std_logic;
signal l3c20_1 : std_logic;
signal l3c19_6 : std_logic;
signal l3c20_2 : std_logic;
signal l3c19_7 : std_logic;
signal l3c20_3 : std_logic;
signal l3c20_4 : std_logic;
signal l3c21_0 : std_logic;
signal l3c20_5 : std_logic;
signal l3c21_1 : std_logic;
signal l3c20_6 : std_logic;
signal l3c21_2 : std_logic;
signal l3c20_7 : std_logic;
signal l3c21_3 : std_logic;
signal l3c20_8 : std_logic;
signal l3c21_4 : std_logic;
signal l3c21_5 : std_logic;
signal l3c22_0 : std_logic;
signal l3c21_6 : std_logic;
signal l3c22_1 : std_logic;
signal l3c21_7 : std_logic;
signal l3c22_2 : std_logic;
signal l3c21_8 : std_logic;
signal l3c22_3 : std_logic;
signal l3c21_9 : std_logic;
signal l3c22_4 : std_logic;
signal l3c22_5 : std_logic;
signal l3c23_0 : std_logic;
signal l3c22_6 : std_logic;
signal l3c23_1 : std_logic;
signal l3c22_7 : std_logic;
signal l3c23_2 : std_logic;
signal l3c22_8 : std_logic;
signal l3c23_3 : std_logic;
signal l3c22_9 : std_logic;
signal l3c23_4 : std_logic;
signal l3c23_5 : std_logic;
signal l3c24_0 : std_logic;
signal l3c23_6 : std_logic;
signal l3c24_1 : std_logic;
signal l3c23_7 : std_logic;
signal l3c24_2 : std_logic;
signal l3c23_8 : std_logic;
signal l3c24_3 : std_logic;
signal l3c23_9 : std_logic;
signal l3c24_4 : std_logic;
signal l3c24_5 : std_logic;
signal l3c25_0 : std_logic;
signal l3c24_6 : std_logic;
signal l3c25_1 : std_logic;
signal l3c24_7 : std_logic;
signal l3c25_2 : std_logic;
signal l3c24_8 : std_logic;
signal l3c25_3 : std_logic;
signal l3c24_9 : std_logic;
signal l3c25_4 : std_logic;
signal l3c25_5 : std_logic;
signal l3c26_0 : std_logic;
signal l3c25_6 : std_logic;
signal l3c26_1 : std_logic;
signal l3c25_7 : std_logic;
signal l3c26_2 : std_logic;
signal l3c25_8 : std_logic;
signal l3c26_3 : std_logic;
signal l3c25_9 : std_logic;
signal l3c26_4 : std_logic;
signal l3c26_5 : std_logic;
signal l3c27_0 : std_logic;
signal l3c26_6 : std_logic;
signal l3c27_1 : std_logic;
signal l3c26_7 : std_logic;
signal l3c27_2 : std_logic;
signal l3c26_8 : std_logic;
signal l3c27_3 : std_logic;
signal l3c26_9 : std_logic;
signal l3c27_4 : std_logic;
signal l3c27_5 : std_logic;
signal l3c28_0 : std_logic;
signal l3c27_6 : std_logic;
signal l3c28_1 : std_logic;
signal l3c27_7 : std_logic;
signal l3c28_2 : std_logic;
signal l3c27_8 : std_logic;
signal l3c28_3 : std_logic;
signal l3c27_9 : std_logic;
signal l3c28_4 : std_logic;
signal l3c28_5 : std_logic;
signal l3c29_0 : std_logic;
signal l3c28_6 : std_logic;
signal l3c29_1 : std_logic;
signal l3c28_7 : std_logic;
signal l3c29_2 : std_logic;
signal l3c28_8 : std_logic;
signal l3c29_3 : std_logic;
signal l3c28_9 : std_logic;
signal l3c29_4 : std_logic;
signal l3c29_5 : std_logic;
signal l3c30_0 : std_logic;
signal l3c29_6 : std_logic;
signal l3c30_1 : std_logic;
signal l3c29_7 : std_logic;
signal l3c30_2 : std_logic;
signal l3c29_8 : std_logic;
signal l3c30_3 : std_logic;
signal l3c30_4 : std_logic;
signal l3c31_0 : std_logic;
signal l3c30_5 : std_logic;
signal l3c31_1 : std_logic;
signal l3c30_6 : std_logic;
signal l3c31_2 : std_logic;
signal l3c30_7 : std_logic;
signal l3c31_3 : std_logic;
signal l3c31_4 : std_logic;
signal l3c32_0 : std_logic;
signal l3c31_5 : std_logic;
signal l3c32_1 : std_logic;
signal l3c31_6 : std_logic;
signal l3c32_2 : std_logic;
signal l3c31_7 : std_logic;
signal l3c32_3 : std_logic;
signal l3c32_4 : std_logic;
signal l3c33_0 : std_logic;
signal l3c32_5 : std_logic;
signal l3c33_1 : std_logic;
signal l3c32_6 : std_logic;
signal l3c33_2 : std_logic;
signal l3c33_3 : std_logic;
signal l3c34_0 : std_logic;
signal l3c33_4 : std_logic;
signal l3c34_1 : std_logic;
signal l3c33_5 : std_logic;
signal l3c34_2 : std_logic;
signal l3c34_3 : std_logic;
signal l3c35_0 : std_logic;
signal l3c34_4 : std_logic;
signal l3c35_1 : std_logic;
signal l3c34_5 : std_logic;
signal l3c35_2 : std_logic;
signal l3c35_3 : std_logic;
signal l3c36_0 : std_logic;
signal l3c35_4 : std_logic;
signal l3c36_1 : std_logic;
signal l3c35_5 : std_logic;
signal l3c36_2 : std_logic;
signal l3c36_3 : std_logic;
signal l3c37_0 : std_logic;
signal l3c36_4 : std_logic;
signal l3c37_1 : std_logic;
signal l3c36_5 : std_logic;
signal l3c37_2 : std_logic;
signal l3c37_3 : std_logic;
signal l3c38_0 : std_logic;
signal l3c37_4 : std_logic;
signal l3c38_1 : std_logic;
signal l3c37_5 : std_logic;
signal l3c38_2 : std_logic;
signal l3c38_3 : std_logic;
signal l3c39_0 : std_logic;
signal l3c38_4 : std_logic;
signal l3c39_1 : std_logic;
signal l3c39_2 : std_logic;
signal l3c40_0 : std_logic;
signal l3c39_3 : std_logic;
signal l3c40_1 : std_logic;
signal l3c40_2 : std_logic;
signal l3c41_0 : std_logic;
signal l3c40_3 : std_logic;
signal l3c41_1 : std_logic;
signal l3c41_2 : std_logic;
signal l3c42_0 : std_logic;
signal l3c42_1 : std_logic;
signal l3c43_0 : std_logic;
signal l3c43_1 : std_logic;
signal l3c44_0 : std_logic;
signal l3c44_1 : std_logic;
signal l3c45_0 : std_logic;
signal l3c45_1 : std_logic;
signal l3c46_0 : std_logic;
signal l3c46_1 : std_logic;
signal l3c47_0 : std_logic;
signal l4c3_0 : std_logic;
signal l4c4_0 : std_logic;
signal l4c4_1 : std_logic;
signal l4c5_0 : std_logic;
signal l4c5_1 : std_logic;
signal l4c6_0 : std_logic;
signal l4c6_1 : std_logic;
signal l4c7_0 : std_logic;
signal l4c7_1 : std_logic;
signal l4c8_0 : std_logic;
signal l4c8_1 : std_logic;
signal l4c9_0 : std_logic;
signal l4c9_1 : std_logic;
signal l4c10_0 : std_logic;
signal l4c9_2 : std_logic;
signal l4c10_1 : std_logic;
signal l4c10_2 : std_logic;
signal l4c11_0 : std_logic;
signal l4c10_3 : std_logic;
signal l4c11_1 : std_logic;
signal l4c11_2 : std_logic;
signal l4c12_0 : std_logic;
signal l4c11_3 : std_logic;
signal l4c12_1 : std_logic;
signal l4c12_2 : std_logic;
signal l4c13_0 : std_logic;
signal l4c12_3 : std_logic;
signal l4c13_1 : std_logic;
signal l4c13_2 : std_logic;
signal l4c14_0 : std_logic;
signal l4c13_3 : std_logic;
signal l4c14_1 : std_logic;
signal l4c14_2 : std_logic;
signal l4c15_0 : std_logic;
signal l4c14_3 : std_logic;
signal l4c15_1 : std_logic;
signal l4c15_2 : std_logic;
signal l4c16_0 : std_logic;
signal l4c15_3 : std_logic;
signal l4c16_1 : std_logic;
signal l4c16_2 : std_logic;
signal l4c17_0 : std_logic;
signal l4c16_3 : std_logic;
signal l4c17_1 : std_logic;
signal l4c16_4 : std_logic;
signal l4c17_2 : std_logic;
signal l4c17_3 : std_logic;
signal l4c18_0 : std_logic;
signal l4c17_4 : std_logic;
signal l4c18_1 : std_logic;
signal l4c17_5 : std_logic;
signal l4c18_2 : std_logic;
signal l4c18_3 : std_logic;
signal l4c19_0 : std_logic;
signal l4c18_4 : std_logic;
signal l4c19_1 : std_logic;
signal l4c18_5 : std_logic;
signal l4c19_2 : std_logic;
signal l4c19_3 : std_logic;
signal l4c20_0 : std_logic;
signal l4c19_4 : std_logic;
signal l4c20_1 : std_logic;
signal l4c19_5 : std_logic;
signal l4c20_2 : std_logic;
signal l4c20_3 : std_logic;
signal l4c21_0 : std_logic;
signal l4c20_4 : std_logic;
signal l4c21_1 : std_logic;
signal l4c20_5 : std_logic;
signal l4c21_2 : std_logic;
signal l4c21_3 : std_logic;
signal l4c22_0 : std_logic;
signal l4c21_4 : std_logic;
signal l4c22_1 : std_logic;
signal l4c21_5 : std_logic;
signal l4c22_2 : std_logic;
signal l4c22_3 : std_logic;
signal l4c23_0 : std_logic;
signal l4c22_4 : std_logic;
signal l4c23_1 : std_logic;
signal l4c22_5 : std_logic;
signal l4c23_2 : std_logic;
signal l4c23_3 : std_logic;
signal l4c24_0 : std_logic;
signal l4c23_4 : std_logic;
signal l4c24_1 : std_logic;
signal l4c23_5 : std_logic;
signal l4c24_2 : std_logic;
signal l4c23_6 : std_logic;
signal l4c24_3 : std_logic;
signal l4c24_4 : std_logic;
signal l4c25_0 : std_logic;
signal l4c24_5 : std_logic;
signal l4c25_1 : std_logic;
signal l4c24_6 : std_logic;
signal l4c25_2 : std_logic;
signal l4c24_7 : std_logic;
signal l4c25_3 : std_logic;
signal l4c25_4 : std_logic;
signal l4c26_0 : std_logic;
signal l4c25_5 : std_logic;
signal l4c26_1 : std_logic;
signal l4c25_6 : std_logic;
signal l4c26_2 : std_logic;
signal l4c25_7 : std_logic;
signal l4c26_3 : std_logic;
signal l4c26_4 : std_logic;
signal l4c27_0 : std_logic;
signal l4c26_5 : std_logic;
signal l4c27_1 : std_logic;
signal l4c26_6 : std_logic;
signal l4c27_2 : std_logic;
signal l4c27_3 : std_logic;
signal l4c28_0 : std_logic;
signal l4c27_4 : std_logic;
signal l4c28_1 : std_logic;
signal l4c27_5 : std_logic;
signal l4c28_2 : std_logic;
signal l4c28_3 : std_logic;
signal l4c29_0 : std_logic;
signal l4c28_4 : std_logic;
signal l4c29_1 : std_logic;
signal l4c28_5 : std_logic;
signal l4c29_2 : std_logic;
signal l4c29_3 : std_logic;
signal l4c30_0 : std_logic;
signal l4c29_4 : std_logic;
signal l4c30_1 : std_logic;
signal l4c29_5 : std_logic;
signal l4c30_2 : std_logic;
signal l4c30_3 : std_logic;
signal l4c31_0 : std_logic;
signal l4c30_4 : std_logic;
signal l4c31_1 : std_logic;
signal l4c30_5 : std_logic;
signal l4c31_2 : std_logic;
signal l4c31_3 : std_logic;
signal l4c32_0 : std_logic;
signal l4c31_4 : std_logic;
signal l4c32_1 : std_logic;
signal l4c31_5 : std_logic;
signal l4c32_2 : std_logic;
signal l4c32_3 : std_logic;
signal l4c33_0 : std_logic;
signal l4c32_4 : std_logic;
signal l4c33_1 : std_logic;
signal l4c32_5 : std_logic;
signal l4c33_2 : std_logic;
signal l4c33_3 : std_logic;
signal l4c34_0 : std_logic;
signal l4c33_4 : std_logic;
signal l4c34_1 : std_logic;
signal l4c34_2 : std_logic;
signal l4c35_0 : std_logic;
signal l4c34_3 : std_logic;
signal l4c35_1 : std_logic;
signal l4c35_2 : std_logic;
signal l4c36_0 : std_logic;
signal l4c35_3 : std_logic;
signal l4c36_1 : std_logic;
signal l4c36_2 : std_logic;
signal l4c37_0 : std_logic;
signal l4c36_3 : std_logic;
signal l4c37_1 : std_logic;
signal l4c37_2 : std_logic;
signal l4c38_0 : std_logic;
signal l4c37_3 : std_logic;
signal l4c38_1 : std_logic;
signal l4c38_2 : std_logic;
signal l4c39_0 : std_logic;
signal l4c38_3 : std_logic;
signal l4c39_1 : std_logic;
signal l4c39_2 : std_logic;
signal l4c40_0 : std_logic;
signal l4c40_1 : std_logic;
signal l4c41_0 : std_logic;
signal l4c41_1 : std_logic;
signal l4c42_0 : std_logic;
signal l4c42_1 : std_logic;
signal l4c43_0 : std_logic;
signal l4c43_1 : std_logic;
signal l4c44_0 : std_logic;
signal l4c44_1 : std_logic;
signal l4c45_0 : std_logic;
signal l4c45_1 : std_logic;
signal l4c46_0 : std_logic;
signal l4c46_1 : std_logic;
signal l4c47_0 : std_logic;
signal l5c4_0 : std_logic;
signal l5c5_0 : std_logic;
signal l5c5_1 : std_logic;
signal l5c6_0 : std_logic;
signal l5c6_1 : std_logic;
signal l5c7_0 : std_logic;
signal l5c7_1 : std_logic;
signal l5c8_0 : std_logic;
signal l5c8_1 : std_logic;
signal l5c9_0 : std_logic;
signal l5c9_1 : std_logic;
signal l5c10_0 : std_logic;
signal l5c10_1 : std_logic;
signal l5c11_0 : std_logic;
signal l5c11_1 : std_logic;
signal l5c12_0 : std_logic;
signal l5c12_1 : std_logic;
signal l5c13_0 : std_logic;
signal l5c13_1 : std_logic;
signal l5c14_0 : std_logic;
signal l5c14_1 : std_logic;
signal l5c15_0 : std_logic;
signal l5c14_2 : std_logic;
signal l5c15_1 : std_logic;
signal l5c15_2 : std_logic;
signal l5c16_0 : std_logic;
signal l5c15_3 : std_logic;
signal l5c16_1 : std_logic;
signal l5c16_2 : std_logic;
signal l5c17_0 : std_logic;
signal l5c16_3 : std_logic;
signal l5c17_1 : std_logic;
signal l5c17_2 : std_logic;
signal l5c18_0 : std_logic;
signal l5c17_3 : std_logic;
signal l5c18_1 : std_logic;
signal l5c18_2 : std_logic;
signal l5c19_0 : std_logic;
signal l5c18_3 : std_logic;
signal l5c19_1 : std_logic;
signal l5c19_2 : std_logic;
signal l5c20_0 : std_logic;
signal l5c19_3 : std_logic;
signal l5c20_1 : std_logic;
signal l5c20_2 : std_logic;
signal l5c21_0 : std_logic;
signal l5c20_3 : std_logic;
signal l5c21_1 : std_logic;
signal l5c21_2 : std_logic;
signal l5c22_0 : std_logic;
signal l5c21_3 : std_logic;
signal l5c22_1 : std_logic;
signal l5c22_2 : std_logic;
signal l5c23_0 : std_logic;
signal l5c22_3 : std_logic;
signal l5c23_1 : std_logic;
signal l5c23_2 : std_logic;
signal l5c24_0 : std_logic;
signal l5c23_3 : std_logic;
signal l5c24_1 : std_logic;
signal l5c24_2 : std_logic;
signal l5c25_0 : std_logic;
signal l5c24_3 : std_logic;
signal l5c25_1 : std_logic;
signal l5c24_4 : std_logic;
signal l5c25_2 : std_logic;
signal l5c25_3 : std_logic;
signal l5c26_0 : std_logic;
signal l5c25_4 : std_logic;
signal l5c26_1 : std_logic;
signal l5c25_5 : std_logic;
signal l5c26_2 : std_logic;
signal l5c26_3 : std_logic;
signal l5c27_0 : std_logic;
signal l5c26_4 : std_logic;
signal l5c27_1 : std_logic;
signal l5c26_5 : std_logic;
signal l5c27_2 : std_logic;
signal l5c27_3 : std_logic;
signal l5c28_0 : std_logic;
signal l5c27_4 : std_logic;
signal l5c28_1 : std_logic;
signal l5c28_2 : std_logic;
signal l5c29_0 : std_logic;
signal l5c28_3 : std_logic;
signal l5c29_1 : std_logic;
signal l5c29_2 : std_logic;
signal l5c30_0 : std_logic;
signal l5c29_3 : std_logic;
signal l5c30_1 : std_logic;
signal l5c30_2 : std_logic;
signal l5c31_0 : std_logic;
signal l5c30_3 : std_logic;
signal l5c31_1 : std_logic;
signal l5c31_2 : std_logic;
signal l5c32_0 : std_logic;
signal l5c31_3 : std_logic;
signal l5c32_1 : std_logic;
signal l5c32_2 : std_logic;
signal l5c33_0 : std_logic;
signal l5c32_3 : std_logic;
signal l5c33_1 : std_logic;
signal l5c33_2 : std_logic;
signal l5c34_0 : std_logic;
signal l5c33_3 : std_logic;
signal l5c34_1 : std_logic;
signal l5c34_2 : std_logic;
signal l5c35_0 : std_logic;
signal l5c34_3 : std_logic;
signal l5c35_1 : std_logic;
signal l5c35_2 : std_logic;
signal l5c36_0 : std_logic;
signal l5c36_1 : std_logic;
signal l5c37_0 : std_logic;
signal l5c37_1 : std_logic;
signal l5c38_0 : std_logic;
signal l5c38_1 : std_logic;
signal l5c39_0 : std_logic;
signal l5c39_1 : std_logic;
signal l5c40_0 : std_logic;
signal l5c40_1 : std_logic;
signal l5c41_0 : std_logic;
signal l5c41_1 : std_logic;
signal l5c42_0 : std_logic;
signal l5c42_1 : std_logic;
signal l5c43_0 : std_logic;
signal l5c43_1 : std_logic;
signal l5c44_0 : std_logic;
signal l5c44_1 : std_logic;
signal l5c45_0 : std_logic;
signal l5c45_1 : std_logic;
signal l5c46_0 : std_logic;
signal l5c46_1 : std_logic;
signal l5c47_0 : std_logic;
signal l5c47_1 : std_logic;
signal l5c48_0 : std_logic;
signal l6c5_0 : std_logic;
signal l6c6_0 : std_logic;
signal l6c6_1 : std_logic;
signal l6c7_0 : std_logic;
signal l6c7_1 : std_logic;
signal l6c8_0 : std_logic;
signal l6c8_1 : std_logic;
signal l6c9_0 : std_logic;
signal l6c9_1 : std_logic;
signal l6c10_0 : std_logic;
signal l6c10_1 : std_logic;
signal l6c11_0 : std_logic;
signal l6c11_1 : std_logic;
signal l6c12_0 : std_logic;
signal l6c12_1 : std_logic;
signal l6c13_0 : std_logic;
signal l6c13_1 : std_logic;
signal l6c14_0 : std_logic;
signal l6c14_1 : std_logic;
signal l6c15_0 : std_logic;
signal l6c15_1 : std_logic;
signal l6c16_0 : std_logic;
signal l6c16_1 : std_logic;
signal l6c17_0 : std_logic;
signal l6c17_1 : std_logic;
signal l6c18_0 : std_logic;
signal l6c18_1 : std_logic;
signal l6c19_0 : std_logic;
signal l6c19_1 : std_logic;
signal l6c20_0 : std_logic;
signal l6c20_1 : std_logic;
signal l6c21_0 : std_logic;
signal l6c21_1 : std_logic;
signal l6c22_0 : std_logic;
signal l6c21_2 : std_logic;
signal l6c22_1 : std_logic;
signal l6c22_2 : std_logic;
signal l6c23_0 : std_logic;
signal l6c22_3 : std_logic;
signal l6c23_1 : std_logic;
signal l6c23_2 : std_logic;
signal l6c24_0 : std_logic;
signal l6c23_3 : std_logic;
signal l6c24_1 : std_logic;
signal l6c24_2 : std_logic;
signal l6c25_0 : std_logic;
signal l6c24_3 : std_logic;
signal l6c25_1 : std_logic;
signal l6c25_2 : std_logic;
signal l6c26_0 : std_logic;
signal l6c25_3 : std_logic;
signal l6c26_1 : std_logic;
signal l6c26_2 : std_logic;
signal l6c27_0 : std_logic;
signal l6c26_3 : std_logic;
signal l6c27_1 : std_logic;
signal l6c27_2 : std_logic;
signal l6c28_0 : std_logic;
signal l6c27_3 : std_logic;
signal l6c28_1 : std_logic;
signal l6c28_2 : std_logic;
signal l6c29_0 : std_logic;
signal l6c28_3 : std_logic;
signal l6c29_1 : std_logic;
signal l6c29_2 : std_logic;
signal l6c30_0 : std_logic;
signal l6c30_1 : std_logic;
signal l6c31_0 : std_logic;
signal l6c31_1 : std_logic;
signal l6c32_0 : std_logic;
signal l6c32_1 : std_logic;
signal l6c33_0 : std_logic;
signal l6c33_1 : std_logic;
signal l6c34_0 : std_logic;
signal l6c34_1 : std_logic;
signal l6c35_0 : std_logic;
signal l6c35_1 : std_logic;
signal l6c36_0 : std_logic;
signal l6c36_1 : std_logic;
signal l6c37_0 : std_logic;
signal l6c37_1 : std_logic;
signal l6c38_0 : std_logic;
signal l6c38_1 : std_logic;
signal l6c39_0 : std_logic;
signal l6c39_1 : std_logic;
signal l6c40_0 : std_logic;
signal l6c40_1 : std_logic;
signal l6c41_0 : std_logic;
signal l6c41_1 : std_logic;
signal l6c42_0 : std_logic;
signal l6c42_1 : std_logic;
signal l6c43_0 : std_logic;
signal l6c43_1 : std_logic;
signal l6c44_0 : std_logic;
signal l6c44_1 : std_logic;
signal l6c45_0 : std_logic;
signal l6c45_1 : std_logic;
signal l6c46_0 : std_logic;
signal l6c46_1 : std_logic;
signal l6c47_0 : std_logic;
signal l6c47_1 : std_logic;
signal l6c48_0 : std_logic;
signal l7c6_0 : std_logic;
signal l7c7_0 : std_logic;
signal l7c7_1 : std_logic;
signal l7c8_0 : std_logic;
signal l7c8_1 : std_logic;
signal l7c9_0 : std_logic;
signal l7c9_1 : std_logic;
signal l7c10_0 : std_logic;
signal l7c10_1 : std_logic;
signal l7c11_0 : std_logic;
signal l7c11_1 : std_logic;
signal l7c12_0 : std_logic;
signal l7c12_1 : std_logic;
signal l7c13_0 : std_logic;
signal l7c13_1 : std_logic;
signal l7c14_0 : std_logic;
signal l7c14_1 : std_logic;
signal l7c15_0 : std_logic;
signal l7c15_1 : std_logic;
signal l7c16_0 : std_logic;
signal l7c16_1 : std_logic;
signal l7c17_0 : std_logic;
signal l7c17_1 : std_logic;
signal l7c18_0 : std_logic;
signal l7c18_1 : std_logic;
signal l7c19_0 : std_logic;
signal l7c19_1 : std_logic;
signal l7c20_0 : std_logic;
signal l7c20_1 : std_logic;
signal l7c21_0 : std_logic;
signal l7c21_1 : std_logic;
signal l7c22_0 : std_logic;
signal l7c22_1 : std_logic;
signal l7c23_0 : std_logic;
signal l7c23_1 : std_logic;
signal l7c24_0 : std_logic;
signal l7c24_1 : std_logic;
signal l7c25_0 : std_logic;
signal l7c25_1 : std_logic;
signal l7c26_0 : std_logic;
signal l7c26_1 : std_logic;
signal l7c27_0 : std_logic;
signal l7c27_1 : std_logic;
signal l7c28_0 : std_logic;
signal l7c28_1 : std_logic;
signal l7c29_0 : std_logic;
signal l7c29_1 : std_logic;
signal l7c30_0 : std_logic;
signal l7c30_1 : std_logic;
signal l7c31_0 : std_logic;
signal l7c31_1 : std_logic;
signal l7c32_0 : std_logic;
signal l7c32_1 : std_logic;
signal l7c33_0 : std_logic;
signal l7c33_1 : std_logic;
signal l7c34_0 : std_logic;
signal l7c34_1 : std_logic;
signal l7c35_0 : std_logic;
signal l7c35_1 : std_logic;
signal l7c36_0 : std_logic;
signal l7c36_1 : std_logic;
signal l7c37_0 : std_logic;
signal l7c37_1 : std_logic;
signal l7c38_0 : std_logic;
signal l7c38_1 : std_logic;
signal l7c39_0 : std_logic;
signal l7c39_1 : std_logic;
signal l7c40_0 : std_logic;
signal l7c40_1 : std_logic;
signal l7c41_0 : std_logic;
signal l7c41_1 : std_logic;
signal l7c42_0 : std_logic;
signal l7c42_1 : std_logic;
signal l7c43_0 : std_logic;
signal l7c43_1 : std_logic;
signal l7c44_0 : std_logic;
signal l7c44_1 : std_logic;
signal l7c45_0 : std_logic;
signal l7c45_1 : std_logic;
signal l7c46_0 : std_logic;
signal l7c46_1 : std_logic;
signal l7c47_0 : std_logic;
signal l7c47_1 : std_logic;
signal l7c48_0 : std_logic;
signal l8c7_0 : std_logic;
signal l8c8_0 : std_logic;
signal l8c8_1 : std_logic;
signal l8c9_0 : std_logic;
signal l8c9_1 : std_logic;
signal l8c10_0 : std_logic;
signal l8c10_1 : std_logic;
signal l8c11_0 : std_logic;
signal l8c11_1 : std_logic;
signal l8c12_0 : std_logic;
signal l8c12_1 : std_logic;
signal l8c13_0 : std_logic;
signal l8c13_1 : std_logic;
signal l8c14_0 : std_logic;
signal l8c14_1 : std_logic;
signal l8c15_0 : std_logic;
signal l8c15_1 : std_logic;
signal l8c16_0 : std_logic;
signal l8c16_1 : std_logic;
signal l8c17_0 : std_logic;
signal l8c17_1 : std_logic;
signal l8c18_0 : std_logic;
signal l8c18_1 : std_logic;
signal l8c19_0 : std_logic;
signal l8c19_1 : std_logic;
signal l8c20_0 : std_logic;
signal l8c20_1 : std_logic;
signal l8c21_0 : std_logic;
signal l8c21_1 : std_logic;
signal l8c22_0 : std_logic;
signal l8c22_1 : std_logic;
signal l8c23_0 : std_logic;
signal l8c23_1 : std_logic;
signal l8c24_0 : std_logic;
signal l8c24_1 : std_logic;
signal l8c25_0 : std_logic;
signal l8c25_1 : std_logic;
signal l8c26_0 : std_logic;
signal l8c26_1 : std_logic;
signal l8c27_0 : std_logic;
signal l8c27_1 : std_logic;
signal l8c28_0 : std_logic;
signal l8c28_1 : std_logic;
signal l8c29_0 : std_logic;
signal l8c29_1 : std_logic;
signal l8c30_0 : std_logic;
signal l8c30_1 : std_logic;
signal l8c31_0 : std_logic;
signal l8c31_1 : std_logic;
signal l8c32_0 : std_logic;
signal l8c32_1 : std_logic;
signal l8c33_0 : std_logic;
signal l8c33_1 : std_logic;
signal l8c34_0 : std_logic;
signal l8c34_1 : std_logic;
signal l8c35_0 : std_logic;
signal l8c35_1 : std_logic;
signal l8c36_0 : std_logic;
signal l8c36_1 : std_logic;
signal l8c37_0 : std_logic;
signal l8c37_1 : std_logic;
signal l8c38_0 : std_logic;
signal l8c38_1 : std_logic;
signal l8c39_0 : std_logic;
signal l8c39_1 : std_logic;
signal l8c40_0 : std_logic;
signal l8c40_1 : std_logic;
signal l8c41_0 : std_logic;
signal l8c41_1 : std_logic;
signal l8c42_0 : std_logic;
signal l8c42_1 : std_logic;
signal l8c43_0 : std_logic;
signal l8c43_1 : std_logic;
signal l8c44_0 : std_logic;
signal l8c44_1 : std_logic;
signal l8c45_0 : std_logic;
signal l8c45_1 : std_logic;
signal l8c46_0 : std_logic;
signal l8c46_1 : std_logic;
signal l8c47_0 : std_logic;
signal l8c47_1 : std_logic;
signal l8c48_0 : std_logic;
signal final_x : std_logic_vector (47 downto 0);
signal final_y : std_logic_vector (47 downto 0);

begin

l1c0_0<= x(0) and y(0);
l1c1_0<= x(1) and y(0);
l1c1_1<= x(0) and y(1);
l1c2_0<= x(2) and y(0);
l1c2_1<= x(1) and y(1);
l1c2_2<= x(0) and y(2);
l1c3_0<= x(3) and y(0);
l1c3_1<= x(2) and y(1);
l1c3_2<= x(1) and y(2);
l1c3_3<= x(0) and y(3);
l1c4_0<= x(4) and y(0);
l1c4_1<= x(3) and y(1);
l1c4_2<= x(2) and y(2);
l1c4_3<= x(1) and y(3);
l1c4_4<= x(0) and y(4);
l1c5_0<= x(5) and y(0);
l1c5_1<= x(4) and y(1);
l1c5_2<= x(3) and y(2);
l1c5_3<= x(2) and y(3);
l1c5_4<= x(1) and y(4);
l1c5_5<= x(0) and y(5);
l1c6_0<= x(6) and y(0);
l1c6_1<= x(5) and y(1);
l1c6_2<= x(4) and y(2);
l1c6_3<= x(3) and y(3);
l1c6_4<= x(2) and y(4);
l1c6_5<= x(1) and y(5);
l1c6_6<= x(0) and y(6);
l1c7_0<= x(7) and y(0);
l1c7_1<= x(6) and y(1);
l1c7_2<= x(5) and y(2);
l1c7_3<= x(4) and y(3);
l1c7_4<= x(3) and y(4);
l1c7_5<= x(2) and y(5);
l1c7_6<= x(1) and y(6);
l1c7_7<= x(0) and y(7);
l1c8_0<= x(8) and y(0);
l1c8_1<= x(7) and y(1);
l1c8_2<= x(6) and y(2);
l1c8_3<= x(5) and y(3);
l1c8_4<= x(4) and y(4);
l1c8_5<= x(3) and y(5);
l1c8_6<= x(2) and y(6);
l1c8_7<= x(1) and y(7);
l1c8_8<= x(0) and y(8);
l1c9_0<= x(9) and y(0);
l1c9_1<= x(8) and y(1);
l1c9_2<= x(7) and y(2);
l1c9_3<= x(6) and y(3);
l1c9_4<= x(5) and y(4);
l1c9_5<= x(4) and y(5);
l1c9_6<= x(3) and y(6);
l1c9_7<= x(2) and y(7);
l1c9_8<= x(1) and y(8);
l1c9_9<= x(0) and y(9);
l1c10_0<= x(10) and y(0);
l1c10_1<= x(9) and y(1);
l1c10_2<= x(8) and y(2);
l1c10_3<= x(7) and y(3);
l1c10_4<= x(6) and y(4);
l1c10_5<= x(5) and y(5);
l1c10_6<= x(4) and y(6);
l1c10_7<= x(3) and y(7);
l1c10_8<= x(2) and y(8);
l1c10_9<= x(1) and y(9);
l1c10_10<= x(0) and y(10);
l1c11_0<= x(11) and y(0);
l1c11_1<= x(10) and y(1);
l1c11_2<= x(9) and y(2);
l1c11_3<= x(8) and y(3);
l1c11_4<= x(7) and y(4);
l1c11_5<= x(6) and y(5);
l1c11_6<= x(5) and y(6);
l1c11_7<= x(4) and y(7);
l1c11_8<= x(3) and y(8);
l1c11_9<= x(2) and y(9);
l1c11_10<= x(1) and y(10);
l1c11_11<= x(0) and y(11);
l1c12_0<= x(12) and y(0);
l1c12_1<= x(11) and y(1);
l1c12_2<= x(10) and y(2);
l1c12_3<= x(9) and y(3);
l1c12_4<= x(8) and y(4);
l1c12_5<= x(7) and y(5);
l1c12_6<= x(6) and y(6);
l1c12_7<= x(5) and y(7);
l1c12_8<= x(4) and y(8);
l1c12_9<= x(3) and y(9);
l1c12_10<= x(2) and y(10);
l1c12_11<= x(1) and y(11);
l1c12_12<= x(0) and y(12);
l1c13_0<= x(13) and y(0);
l1c13_1<= x(12) and y(1);
l1c13_2<= x(11) and y(2);
l1c13_3<= x(10) and y(3);
l1c13_4<= x(9) and y(4);
l1c13_5<= x(8) and y(5);
l1c13_6<= x(7) and y(6);
l1c13_7<= x(6) and y(7);
l1c13_8<= x(5) and y(8);
l1c13_9<= x(4) and y(9);
l1c13_10<= x(3) and y(10);
l1c13_11<= x(2) and y(11);
l1c13_12<= x(1) and y(12);
l1c13_13<= x(0) and y(13);
l1c14_0<= x(14) and y(0);
l1c14_1<= x(13) and y(1);
l1c14_2<= x(12) and y(2);
l1c14_3<= x(11) and y(3);
l1c14_4<= x(10) and y(4);
l1c14_5<= x(9) and y(5);
l1c14_6<= x(8) and y(6);
l1c14_7<= x(7) and y(7);
l1c14_8<= x(6) and y(8);
l1c14_9<= x(5) and y(9);
l1c14_10<= x(4) and y(10);
l1c14_11<= x(3) and y(11);
l1c14_12<= x(2) and y(12);
l1c14_13<= x(1) and y(13);
l1c14_14<= x(0) and y(14);
l1c15_0<= x(15) and y(0);
l1c15_1<= x(14) and y(1);
l1c15_2<= x(13) and y(2);
l1c15_3<= x(12) and y(3);
l1c15_4<= x(11) and y(4);
l1c15_5<= x(10) and y(5);
l1c15_6<= x(9) and y(6);
l1c15_7<= x(8) and y(7);
l1c15_8<= x(7) and y(8);
l1c15_9<= x(6) and y(9);
l1c15_10<= x(5) and y(10);
l1c15_11<= x(4) and y(11);
l1c15_12<= x(3) and y(12);
l1c15_13<= x(2) and y(13);
l1c15_14<= x(1) and y(14);
l1c15_15<= x(0) and y(15);
l1c16_0<= x(16) and y(0);
l1c16_1<= x(15) and y(1);
l1c16_2<= x(14) and y(2);
l1c16_3<= x(13) and y(3);
l1c16_4<= x(12) and y(4);
l1c16_5<= x(11) and y(5);
l1c16_6<= x(10) and y(6);
l1c16_7<= x(9) and y(7);
l1c16_8<= x(8) and y(8);
l1c16_9<= x(7) and y(9);
l1c16_10<= x(6) and y(10);
l1c16_11<= x(5) and y(11);
l1c16_12<= x(4) and y(12);
l1c16_13<= x(3) and y(13);
l1c16_14<= x(2) and y(14);
l1c16_15<= x(1) and y(15);
l1c16_16<= x(0) and y(16);
l1c17_0<= x(17) and y(0);
l1c17_1<= x(16) and y(1);
l1c17_2<= x(15) and y(2);
l1c17_3<= x(14) and y(3);
l1c17_4<= x(13) and y(4);
l1c17_5<= x(12) and y(5);
l1c17_6<= x(11) and y(6);
l1c17_7<= x(10) and y(7);
l1c17_8<= x(9) and y(8);
l1c17_9<= x(8) and y(9);
l1c17_10<= x(7) and y(10);
l1c17_11<= x(6) and y(11);
l1c17_12<= x(5) and y(12);
l1c17_13<= x(4) and y(13);
l1c17_14<= x(3) and y(14);
l1c17_15<= x(2) and y(15);
l1c17_16<= x(1) and y(16);
l1c17_17<= x(0) and y(17);
l1c18_0<= x(18) and y(0);
l1c18_1<= x(17) and y(1);
l1c18_2<= x(16) and y(2);
l1c18_3<= x(15) and y(3);
l1c18_4<= x(14) and y(4);
l1c18_5<= x(13) and y(5);
l1c18_6<= x(12) and y(6);
l1c18_7<= x(11) and y(7);
l1c18_8<= x(10) and y(8);
l1c18_9<= x(9) and y(9);
l1c18_10<= x(8) and y(10);
l1c18_11<= x(7) and y(11);
l1c18_12<= x(6) and y(12);
l1c18_13<= x(5) and y(13);
l1c18_14<= x(4) and y(14);
l1c18_15<= x(3) and y(15);
l1c18_16<= x(2) and y(16);
l1c18_17<= x(1) and y(17);
l1c18_18<= x(0) and y(18);
l1c19_0<= x(19) and y(0);
l1c19_1<= x(18) and y(1);
l1c19_2<= x(17) and y(2);
l1c19_3<= x(16) and y(3);
l1c19_4<= x(15) and y(4);
l1c19_5<= x(14) and y(5);
l1c19_6<= x(13) and y(6);
l1c19_7<= x(12) and y(7);
l1c19_8<= x(11) and y(8);
l1c19_9<= x(10) and y(9);
l1c19_10<= x(9) and y(10);
l1c19_11<= x(8) and y(11);
l1c19_12<= x(7) and y(12);
l1c19_13<= x(6) and y(13);
l1c19_14<= x(5) and y(14);
l1c19_15<= x(4) and y(15);
l1c19_16<= x(3) and y(16);
l1c19_17<= x(2) and y(17);
l1c19_18<= x(1) and y(18);
l1c19_19<= x(0) and y(19);
l1c20_0<= x(20) and y(0);
l1c20_1<= x(19) and y(1);
l1c20_2<= x(18) and y(2);
l1c20_3<= x(17) and y(3);
l1c20_4<= x(16) and y(4);
l1c20_5<= x(15) and y(5);
l1c20_6<= x(14) and y(6);
l1c20_7<= x(13) and y(7);
l1c20_8<= x(12) and y(8);
l1c20_9<= x(11) and y(9);
l1c20_10<= x(10) and y(10);
l1c20_11<= x(9) and y(11);
l1c20_12<= x(8) and y(12);
l1c20_13<= x(7) and y(13);
l1c20_14<= x(6) and y(14);
l1c20_15<= x(5) and y(15);
l1c20_16<= x(4) and y(16);
l1c20_17<= x(3) and y(17);
l1c20_18<= x(2) and y(18);
l1c20_19<= x(1) and y(19);
l1c20_20<= x(0) and y(20);
l1c21_0<= x(21) and y(0);
l1c21_1<= x(20) and y(1);
l1c21_2<= x(19) and y(2);
l1c21_3<= x(18) and y(3);
l1c21_4<= x(17) and y(4);
l1c21_5<= x(16) and y(5);
l1c21_6<= x(15) and y(6);
l1c21_7<= x(14) and y(7);
l1c21_8<= x(13) and y(8);
l1c21_9<= x(12) and y(9);
l1c21_10<= x(11) and y(10);
l1c21_11<= x(10) and y(11);
l1c21_12<= x(9) and y(12);
l1c21_13<= x(8) and y(13);
l1c21_14<= x(7) and y(14);
l1c21_15<= x(6) and y(15);
l1c21_16<= x(5) and y(16);
l1c21_17<= x(4) and y(17);
l1c21_18<= x(3) and y(18);
l1c21_19<= x(2) and y(19);
l1c21_20<= x(1) and y(20);
l1c21_21<= x(0) and y(21);
l1c22_0<= x(22) and y(0);
l1c22_1<= x(21) and y(1);
l1c22_2<= x(20) and y(2);
l1c22_3<= x(19) and y(3);
l1c22_4<= x(18) and y(4);
l1c22_5<= x(17) and y(5);
l1c22_6<= x(16) and y(6);
l1c22_7<= x(15) and y(7);
l1c22_8<= x(14) and y(8);
l1c22_9<= x(13) and y(9);
l1c22_10<= x(12) and y(10);
l1c22_11<= x(11) and y(11);
l1c22_12<= x(10) and y(12);
l1c22_13<= x(9) and y(13);
l1c22_14<= x(8) and y(14);
l1c22_15<= x(7) and y(15);
l1c22_16<= x(6) and y(16);
l1c22_17<= x(5) and y(17);
l1c22_18<= x(4) and y(18);
l1c22_19<= x(3) and y(19);
l1c22_20<= x(2) and y(20);
l1c22_21<= x(1) and y(21);
l1c22_22<= x(0) and y(22);
l1c23_0<= x(23) and y(0);
l1c23_1<= x(22) and y(1);
l1c23_2<= x(21) and y(2);
l1c23_3<= x(20) and y(3);
l1c23_4<= x(19) and y(4);
l1c23_5<= x(18) and y(5);
l1c23_6<= x(17) and y(6);
l1c23_7<= x(16) and y(7);
l1c23_8<= x(15) and y(8);
l1c23_9<= x(14) and y(9);
l1c23_10<= x(13) and y(10);
l1c23_11<= x(12) and y(11);
l1c23_12<= x(11) and y(12);
l1c23_13<= x(10) and y(13);
l1c23_14<= x(9) and y(14);
l1c23_15<= x(8) and y(15);
l1c23_16<= x(7) and y(16);
l1c23_17<= x(6) and y(17);
l1c23_18<= x(5) and y(18);
l1c23_19<= x(4) and y(19);
l1c23_20<= x(3) and y(20);
l1c23_21<= x(2) and y(21);
l1c23_22<= x(1) and y(22);
l1c23_23<= x(0) and y(23);
l1c24_0<= x(23) and y(1);
l1c24_1<= x(22) and y(2);
l1c24_2<= x(21) and y(3);
l1c24_3<= x(20) and y(4);
l1c24_4<= x(19) and y(5);
l1c24_5<= x(18) and y(6);
l1c24_6<= x(17) and y(7);
l1c24_7<= x(16) and y(8);
l1c24_8<= x(15) and y(9);
l1c24_9<= x(14) and y(10);
l1c24_10<= x(13) and y(11);
l1c24_11<= x(12) and y(12);
l1c24_12<= x(11) and y(13);
l1c24_13<= x(10) and y(14);
l1c24_14<= x(9) and y(15);
l1c24_15<= x(8) and y(16);
l1c24_16<= x(7) and y(17);
l1c24_17<= x(6) and y(18);
l1c24_18<= x(5) and y(19);
l1c24_19<= x(4) and y(20);
l1c24_20<= x(3) and y(21);
l1c24_21<= x(2) and y(22);
l1c24_22<= x(1) and y(23);
l1c25_0<= x(23) and y(2);
l1c25_1<= x(22) and y(3);
l1c25_2<= x(21) and y(4);
l1c25_3<= x(20) and y(5);
l1c25_4<= x(19) and y(6);
l1c25_5<= x(18) and y(7);
l1c25_6<= x(17) and y(8);
l1c25_7<= x(16) and y(9);
l1c25_8<= x(15) and y(10);
l1c25_9<= x(14) and y(11);
l1c25_10<= x(13) and y(12);
l1c25_11<= x(12) and y(13);
l1c25_12<= x(11) and y(14);
l1c25_13<= x(10) and y(15);
l1c25_14<= x(9) and y(16);
l1c25_15<= x(8) and y(17);
l1c25_16<= x(7) and y(18);
l1c25_17<= x(6) and y(19);
l1c25_18<= x(5) and y(20);
l1c25_19<= x(4) and y(21);
l1c25_20<= x(3) and y(22);
l1c25_21<= x(2) and y(23);
l1c26_0<= x(23) and y(3);
l1c26_1<= x(22) and y(4);
l1c26_2<= x(21) and y(5);
l1c26_3<= x(20) and y(6);
l1c26_4<= x(19) and y(7);
l1c26_5<= x(18) and y(8);
l1c26_6<= x(17) and y(9);
l1c26_7<= x(16) and y(10);
l1c26_8<= x(15) and y(11);
l1c26_9<= x(14) and y(12);
l1c26_10<= x(13) and y(13);
l1c26_11<= x(12) and y(14);
l1c26_12<= x(11) and y(15);
l1c26_13<= x(10) and y(16);
l1c26_14<= x(9) and y(17);
l1c26_15<= x(8) and y(18);
l1c26_16<= x(7) and y(19);
l1c26_17<= x(6) and y(20);
l1c26_18<= x(5) and y(21);
l1c26_19<= x(4) and y(22);
l1c26_20<= x(3) and y(23);
l1c27_0<= x(23) and y(4);
l1c27_1<= x(22) and y(5);
l1c27_2<= x(21) and y(6);
l1c27_3<= x(20) and y(7);
l1c27_4<= x(19) and y(8);
l1c27_5<= x(18) and y(9);
l1c27_6<= x(17) and y(10);
l1c27_7<= x(16) and y(11);
l1c27_8<= x(15) and y(12);
l1c27_9<= x(14) and y(13);
l1c27_10<= x(13) and y(14);
l1c27_11<= x(12) and y(15);
l1c27_12<= x(11) and y(16);
l1c27_13<= x(10) and y(17);
l1c27_14<= x(9) and y(18);
l1c27_15<= x(8) and y(19);
l1c27_16<= x(7) and y(20);
l1c27_17<= x(6) and y(21);
l1c27_18<= x(5) and y(22);
l1c27_19<= x(4) and y(23);
l1c28_0<= x(23) and y(5);
l1c28_1<= x(22) and y(6);
l1c28_2<= x(21) and y(7);
l1c28_3<= x(20) and y(8);
l1c28_4<= x(19) and y(9);
l1c28_5<= x(18) and y(10);
l1c28_6<= x(17) and y(11);
l1c28_7<= x(16) and y(12);
l1c28_8<= x(15) and y(13);
l1c28_9<= x(14) and y(14);
l1c28_10<= x(13) and y(15);
l1c28_11<= x(12) and y(16);
l1c28_12<= x(11) and y(17);
l1c28_13<= x(10) and y(18);
l1c28_14<= x(9) and y(19);
l1c28_15<= x(8) and y(20);
l1c28_16<= x(7) and y(21);
l1c28_17<= x(6) and y(22);
l1c28_18<= x(5) and y(23);
l1c29_0<= x(23) and y(6);
l1c29_1<= x(22) and y(7);
l1c29_2<= x(21) and y(8);
l1c29_3<= x(20) and y(9);
l1c29_4<= x(19) and y(10);
l1c29_5<= x(18) and y(11);
l1c29_6<= x(17) and y(12);
l1c29_7<= x(16) and y(13);
l1c29_8<= x(15) and y(14);
l1c29_9<= x(14) and y(15);
l1c29_10<= x(13) and y(16);
l1c29_11<= x(12) and y(17);
l1c29_12<= x(11) and y(18);
l1c29_13<= x(10) and y(19);
l1c29_14<= x(9) and y(20);
l1c29_15<= x(8) and y(21);
l1c29_16<= x(7) and y(22);
l1c29_17<= x(6) and y(23);
l1c30_0<= x(23) and y(7);
l1c30_1<= x(22) and y(8);
l1c30_2<= x(21) and y(9);
l1c30_3<= x(20) and y(10);
l1c30_4<= x(19) and y(11);
l1c30_5<= x(18) and y(12);
l1c30_6<= x(17) and y(13);
l1c30_7<= x(16) and y(14);
l1c30_8<= x(15) and y(15);
l1c30_9<= x(14) and y(16);
l1c30_10<= x(13) and y(17);
l1c30_11<= x(12) and y(18);
l1c30_12<= x(11) and y(19);
l1c30_13<= x(10) and y(20);
l1c30_14<= x(9) and y(21);
l1c30_15<= x(8) and y(22);
l1c30_16<= x(7) and y(23);
l1c31_0<= x(23) and y(8);
l1c31_1<= x(22) and y(9);
l1c31_2<= x(21) and y(10);
l1c31_3<= x(20) and y(11);
l1c31_4<= x(19) and y(12);
l1c31_5<= x(18) and y(13);
l1c31_6<= x(17) and y(14);
l1c31_7<= x(16) and y(15);
l1c31_8<= x(15) and y(16);
l1c31_9<= x(14) and y(17);
l1c31_10<= x(13) and y(18);
l1c31_11<= x(12) and y(19);
l1c31_12<= x(11) and y(20);
l1c31_13<= x(10) and y(21);
l1c31_14<= x(9) and y(22);
l1c31_15<= x(8) and y(23);
l1c32_0<= x(23) and y(9);
l1c32_1<= x(22) and y(10);
l1c32_2<= x(21) and y(11);
l1c32_3<= x(20) and y(12);
l1c32_4<= x(19) and y(13);
l1c32_5<= x(18) and y(14);
l1c32_6<= x(17) and y(15);
l1c32_7<= x(16) and y(16);
l1c32_8<= x(15) and y(17);
l1c32_9<= x(14) and y(18);
l1c32_10<= x(13) and y(19);
l1c32_11<= x(12) and y(20);
l1c32_12<= x(11) and y(21);
l1c32_13<= x(10) and y(22);
l1c32_14<= x(9) and y(23);
l1c33_0<= x(23) and y(10);
l1c33_1<= x(22) and y(11);
l1c33_2<= x(21) and y(12);
l1c33_3<= x(20) and y(13);
l1c33_4<= x(19) and y(14);
l1c33_5<= x(18) and y(15);
l1c33_6<= x(17) and y(16);
l1c33_7<= x(16) and y(17);
l1c33_8<= x(15) and y(18);
l1c33_9<= x(14) and y(19);
l1c33_10<= x(13) and y(20);
l1c33_11<= x(12) and y(21);
l1c33_12<= x(11) and y(22);
l1c33_13<= x(10) and y(23);
l1c34_0<= x(23) and y(11);
l1c34_1<= x(22) and y(12);
l1c34_2<= x(21) and y(13);
l1c34_3<= x(20) and y(14);
l1c34_4<= x(19) and y(15);
l1c34_5<= x(18) and y(16);
l1c34_6<= x(17) and y(17);
l1c34_7<= x(16) and y(18);
l1c34_8<= x(15) and y(19);
l1c34_9<= x(14) and y(20);
l1c34_10<= x(13) and y(21);
l1c34_11<= x(12) and y(22);
l1c34_12<= x(11) and y(23);
l1c35_0<= x(23) and y(12);
l1c35_1<= x(22) and y(13);
l1c35_2<= x(21) and y(14);
l1c35_3<= x(20) and y(15);
l1c35_4<= x(19) and y(16);
l1c35_5<= x(18) and y(17);
l1c35_6<= x(17) and y(18);
l1c35_7<= x(16) and y(19);
l1c35_8<= x(15) and y(20);
l1c35_9<= x(14) and y(21);
l1c35_10<= x(13) and y(22);
l1c35_11<= x(12) and y(23);
l1c36_0<= x(23) and y(13);
l1c36_1<= x(22) and y(14);
l1c36_2<= x(21) and y(15);
l1c36_3<= x(20) and y(16);
l1c36_4<= x(19) and y(17);
l1c36_5<= x(18) and y(18);
l1c36_6<= x(17) and y(19);
l1c36_7<= x(16) and y(20);
l1c36_8<= x(15) and y(21);
l1c36_9<= x(14) and y(22);
l1c36_10<= x(13) and y(23);
l1c37_0<= x(23) and y(14);
l1c37_1<= x(22) and y(15);
l1c37_2<= x(21) and y(16);
l1c37_3<= x(20) and y(17);
l1c37_4<= x(19) and y(18);
l1c37_5<= x(18) and y(19);
l1c37_6<= x(17) and y(20);
l1c37_7<= x(16) and y(21);
l1c37_8<= x(15) and y(22);
l1c37_9<= x(14) and y(23);
l1c38_0<= x(23) and y(15);
l1c38_1<= x(22) and y(16);
l1c38_2<= x(21) and y(17);
l1c38_3<= x(20) and y(18);
l1c38_4<= x(19) and y(19);
l1c38_5<= x(18) and y(20);
l1c38_6<= x(17) and y(21);
l1c38_7<= x(16) and y(22);
l1c38_8<= x(15) and y(23);
l1c39_0<= x(23) and y(16);
l1c39_1<= x(22) and y(17);
l1c39_2<= x(21) and y(18);
l1c39_3<= x(20) and y(19);
l1c39_4<= x(19) and y(20);
l1c39_5<= x(18) and y(21);
l1c39_6<= x(17) and y(22);
l1c39_7<= x(16) and y(23);
l1c40_0<= x(23) and y(17);
l1c40_1<= x(22) and y(18);
l1c40_2<= x(21) and y(19);
l1c40_3<= x(20) and y(20);
l1c40_4<= x(19) and y(21);
l1c40_5<= x(18) and y(22);
l1c40_6<= x(17) and y(23);
l1c41_0<= x(23) and y(18);
l1c41_1<= x(22) and y(19);
l1c41_2<= x(21) and y(20);
l1c41_3<= x(20) and y(21);
l1c41_4<= x(19) and y(22);
l1c41_5<= x(18) and y(23);
l1c42_0<= x(23) and y(19);
l1c42_1<= x(22) and y(20);
l1c42_2<= x(21) and y(21);
l1c42_3<= x(20) and y(22);
l1c42_4<= x(19) and y(23);
l1c43_0<= x(23) and y(20);
l1c43_1<= x(22) and y(21);
l1c43_2<= x(21) and y(22);
l1c43_3<= x(20) and y(23);
l1c44_0<= x(23) and y(21);
l1c44_1<= x(22) and y(22);
l1c44_2<= x(21) and y(23);
l1c45_0<= x(23) and y(22);
l1c45_1<= x(22) and y(23);
l1c46_0<= x(23) and y(23);

halfadder0: half_adder port map(x => l1c1_0, y => l1c1_1, s => l2c1_0, cout => l2c2_0);
halfadder1: half_adder port map(x => l1c4_3, y => l1c4_4, s => l2c4_2, cout => l2c5_1);
halfadder2: half_adder port map(x => l1c7_6, y => l1c7_7, s => l2c7_4, cout => l2c8_2);
halfadder3: half_adder port map(x => l1c10_9, y => l1c10_10, s => l2c10_6, cout => l2c11_3);
halfadder4: half_adder port map(x => l1c13_12, y => l1c13_13, s => l2c13_8, cout => l2c14_4);
halfadder5: half_adder port map(x => l1c16_15, y => l1c16_16, s => l2c16_10, cout => l2c17_5);
halfadder6: half_adder port map(x => l1c19_18, y => l1c19_19, s => l2c19_12, cout => l2c20_6);
halfadder7: half_adder port map(x => l1c22_21, y => l1c22_22, s => l2c22_14, cout => l2c23_7);
halfadder8: half_adder port map(x => l1c24_21, y => l1c24_22, s => l2c24_15, cout => l2c25_7);
halfadder9: half_adder port map(x => l1c27_18, y => l1c27_19, s => l2c27_13, cout => l2c28_6);
halfadder10: half_adder port map(x => l1c30_15, y => l1c30_16, s => l2c30_11, cout => l2c31_5);
halfadder11: half_adder port map(x => l1c33_12, y => l1c33_13, s => l2c33_9, cout => l2c34_4);
halfadder12: half_adder port map(x => l1c36_9, y => l1c36_10, s => l2c36_7, cout => l2c37_3);
halfadder13: half_adder port map(x => l1c39_6, y => l1c39_7, s => l2c39_5, cout => l2c40_2);
halfadder14: half_adder port map(x => l1c42_3, y => l1c42_4, s => l2c42_3, cout => l2c43_1);
halfadder15: half_adder port map(x => l1c45_0, y => l1c45_1, s => l2c45_1, cout => l2c46_0);
halfadder16: half_adder port map(x => l2c2_0, y => l2c2_1, s => l3c2_0, cout => l3c3_0);
halfadder17: half_adder port map(x => l2c6_3, y => l1c6_6, s => l3c6_2, cout => l3c7_1);
halfadder18: half_adder port map(x => l2c7_3, y => l2c7_4, s => l3c7_3, cout => l3c8_1);
halfadder19: half_adder port map(x => l2c11_6, y => l2c11_7, s => l3c11_4, cout => l3c12_2);
halfadder20: half_adder port map(x => l2c15_9, y => l1c15_15, s => l3c15_6, cout => l3c16_3);
halfadder21: half_adder port map(x => l2c16_9, y => l2c16_10, s => l3c16_7, cout => l3c17_3);
halfadder22: half_adder port map(x => l2c20_12, y => l2c20_13, s => l3c20_8, cout => l3c21_4);
halfadder23: half_adder port map(x => l2c26_12, y => l2c26_13, s => l3c26_9, cout => l3c27_4);
halfadder24: half_adder port map(x => l2c27_12, y => l2c27_13, s => l3c27_9, cout => l3c28_4);
halfadder25: half_adder port map(x => l2c28_12, y => l1c28_18, s => l3c28_9, cout => l3c29_4);
halfadder26: half_adder port map(x => l2c35_6, y => l2c35_7, s => l3c35_5, cout => l3c36_2);
halfadder27: half_adder port map(x => l2c36_6, y => l2c36_7, s => l3c36_5, cout => l3c37_2);
halfadder28: half_adder port map(x => l2c37_6, y => l1c37_9, s => l3c37_5, cout => l3c38_2);
halfadder29: half_adder port map(x => l2c44_0, y => l2c44_1, s => l3c44_1, cout => l3c45_0);
halfadder30: half_adder port map(x => l2c45_0, y => l2c45_1, s => l3c45_1, cout => l3c46_0);
halfadder31: half_adder port map(x => l2c46_0, y => l1c46_0, s => l3c46_1, cout => l3c47_0);
halfadder32: half_adder port map(x => l3c3_0, y => l3c3_1, s => l4c3_0, cout => l4c4_0);
halfadder33: half_adder port map(x => l3c4_0, y => l3c4_1, s => l4c4_1, cout => l4c5_0);
halfadder34: half_adder port map(x => l3c9_3, y => l1c9_9, s => l4c9_2, cout => l4c10_1);
halfadder35: half_adder port map(x => l3c10_3, y => l2c10_6, s => l4c10_3, cout => l4c11_1);
halfadder36: half_adder port map(x => l3c11_3, y => l3c11_4, s => l4c11_3, cout => l4c12_1);
halfadder37: half_adder port map(x => l3c16_6, y => l3c16_7, s => l4c16_4, cout => l4c17_2);
halfadder38: half_adder port map(x => l3c17_6, y => l3c17_7, s => l4c17_5, cout => l4c18_2);
halfadder39: half_adder port map(x => l3c23_9, y => l2c23_15, s => l4c23_6, cout => l4c24_3);
halfadder40: half_adder port map(x => l3c24_9, y => l2c24_15, s => l4c24_7, cout => l4c25_3);
halfadder41: half_adder port map(x => l3c25_9, y => l1c25_21, s => l4c25_7, cout => l4c26_3);
halfadder42: half_adder port map(x => l3c30_6, y => l3c30_7, s => l4c30_5, cout => l4c31_2);
halfadder43: half_adder port map(x => l3c31_6, y => l3c31_7, s => l4c31_5, cout => l4c32_2);
halfadder44: half_adder port map(x => l3c32_6, y => l2c32_9, s => l4c32_5, cout => l4c33_2);
halfadder45: half_adder port map(x => l3c38_3, y => l3c38_4, s => l4c38_3, cout => l4c39_1);
halfadder46: half_adder port map(x => l3c44_0, y => l3c44_1, s => l4c44_1, cout => l4c45_0);
halfadder47: half_adder port map(x => l3c45_0, y => l3c45_1, s => l4c45_1, cout => l4c46_0);
halfadder48: half_adder port map(x => l3c46_0, y => l3c46_1, s => l4c46_1, cout => l4c47_0);
halfadder49: half_adder port map(x => l4c4_0, y => l4c4_1, s => l5c4_0, cout => l5c5_0);
halfadder50: half_adder port map(x => l4c5_0, y => l4c5_1, s => l5c5_1, cout => l5c6_0);
halfadder51: half_adder port map(x => l4c6_0, y => l4c6_1, s => l5c6_1, cout => l5c7_0);
halfadder52: half_adder port map(x => l4c14_3, y => l2c14_9, s => l5c14_2, cout => l5c15_1);
halfadder53: half_adder port map(x => l4c15_3, y => l3c15_6, s => l5c15_3, cout => l5c16_1);
halfadder54: half_adder port map(x => l4c16_3, y => l4c16_4, s => l5c16_3, cout => l5c17_1);
halfadder55: half_adder port map(x => l4c24_6, y => l4c24_7, s => l5c24_4, cout => l5c25_2);
halfadder56: half_adder port map(x => l4c25_6, y => l4c25_7, s => l5c25_5, cout => l5c26_2);
halfadder57: half_adder port map(x => l4c26_6, y => l3c26_9, s => l5c26_5, cout => l5c27_2);
halfadder58: half_adder port map(x => l4c34_3, y => l1c34_12, s => l5c34_3, cout => l5c35_1);
halfadder59: half_adder port map(x => l4c42_0, y => l4c42_1, s => l5c42_1, cout => l5c43_0);
halfadder60: half_adder port map(x => l4c43_0, y => l4c43_1, s => l5c43_1, cout => l5c44_0);
halfadder61: half_adder port map(x => l4c44_0, y => l4c44_1, s => l5c44_1, cout => l5c45_0);
halfadder62: half_adder port map(x => l4c45_0, y => l4c45_1, s => l5c45_1, cout => l5c46_0);
halfadder63: half_adder port map(x => l4c46_0, y => l4c46_1, s => l5c46_1, cout => l5c47_0);
halfadder64: half_adder port map(x => l4c47_0, y => l3c47_0, s => l5c47_1, cout => l5c48_0);
halfadder65: half_adder port map(x => l5c5_0, y => l5c5_1, s => l6c5_0, cout => l6c6_0);
halfadder66: half_adder port map(x => l5c6_0, y => l5c6_1, s => l6c6_1, cout => l6c7_0);
halfadder67: half_adder port map(x => l5c7_0, y => l5c7_1, s => l6c7_1, cout => l6c8_0);
halfadder68: half_adder port map(x => l5c8_0, y => l5c8_1, s => l6c8_1, cout => l6c9_0);
halfadder69: half_adder port map(x => l5c9_0, y => l5c9_1, s => l6c9_1, cout => l6c10_0);
halfadder70: half_adder port map(x => l5c21_3, y => l3c21_9, s => l6c21_2, cout => l6c22_1);
halfadder71: half_adder port map(x => l5c22_3, y => l3c22_9, s => l6c22_3, cout => l6c23_1);
halfadder72: half_adder port map(x => l5c23_3, y => l4c23_6, s => l6c23_3, cout => l6c24_1);
halfadder73: half_adder port map(x => l5c24_3, y => l5c24_4, s => l6c24_3, cout => l6c25_1);
halfadder74: half_adder port map(x => l5c28_3, y => l3c28_9, s => l6c28_3, cout => l6c29_1);
halfadder75: half_adder port map(x => l5c40_0, y => l5c40_1, s => l6c40_1, cout => l6c41_0);
halfadder76: half_adder port map(x => l5c41_0, y => l5c41_1, s => l6c41_1, cout => l6c42_0);
halfadder77: half_adder port map(x => l5c42_0, y => l5c42_1, s => l6c42_1, cout => l6c43_0);
halfadder78: half_adder port map(x => l5c43_0, y => l5c43_1, s => l6c43_1, cout => l6c44_0);
halfadder79: half_adder port map(x => l5c44_0, y => l5c44_1, s => l6c44_1, cout => l6c45_0);
halfadder80: half_adder port map(x => l5c45_0, y => l5c45_1, s => l6c45_1, cout => l6c46_0);
halfadder81: half_adder port map(x => l5c46_0, y => l5c46_1, s => l6c46_1, cout => l6c47_0);
halfadder82: half_adder port map(x => l5c47_0, y => l5c47_1, s => l6c47_1, cout => l6c48_0);
halfadder83: half_adder port map(x => l6c6_0, y => l6c6_1, s => l7c6_0, cout => l7c7_0);
halfadder84: half_adder port map(x => l6c7_0, y => l6c7_1, s => l7c7_1, cout => l7c8_0);
halfadder85: half_adder port map(x => l6c8_0, y => l6c8_1, s => l7c8_1, cout => l7c9_0);
halfadder86: half_adder port map(x => l6c9_0, y => l6c9_1, s => l7c9_1, cout => l7c10_0);
halfadder87: half_adder port map(x => l6c10_0, y => l6c10_1, s => l7c10_1, cout => l7c11_0);
halfadder88: half_adder port map(x => l6c11_0, y => l6c11_1, s => l7c11_1, cout => l7c12_0);
halfadder89: half_adder port map(x => l6c12_0, y => l6c12_1, s => l7c12_1, cout => l7c13_0);
halfadder90: half_adder port map(x => l6c13_0, y => l6c13_1, s => l7c13_1, cout => l7c14_0);
halfadder91: half_adder port map(x => l6c14_0, y => l6c14_1, s => l7c14_1, cout => l7c15_0);
halfadder92: half_adder port map(x => l6c36_0, y => l6c36_1, s => l7c36_1, cout => l7c37_0);
halfadder93: half_adder port map(x => l6c37_0, y => l6c37_1, s => l7c37_1, cout => l7c38_0);
halfadder94: half_adder port map(x => l6c38_0, y => l6c38_1, s => l7c38_1, cout => l7c39_0);
halfadder95: half_adder port map(x => l6c39_0, y => l6c39_1, s => l7c39_1, cout => l7c40_0);
halfadder96: half_adder port map(x => l6c40_0, y => l6c40_1, s => l7c40_1, cout => l7c41_0);
halfadder97: half_adder port map(x => l6c41_0, y => l6c41_1, s => l7c41_1, cout => l7c42_0);
halfadder98: half_adder port map(x => l6c42_0, y => l6c42_1, s => l7c42_1, cout => l7c43_0);
halfadder99: half_adder port map(x => l6c43_0, y => l6c43_1, s => l7c43_1, cout => l7c44_0);
halfadder100: half_adder port map(x => l6c44_0, y => l6c44_1, s => l7c44_1, cout => l7c45_0);
halfadder101: half_adder port map(x => l6c45_0, y => l6c45_1, s => l7c45_1, cout => l7c46_0);
halfadder102: half_adder port map(x => l6c46_0, y => l6c46_1, s => l7c46_1, cout => l7c47_0);
halfadder103: half_adder port map(x => l6c47_0, y => l6c47_1, s => l7c47_1, cout => l7c48_0);
halfadder104: half_adder port map(x => l7c7_0, y => l7c7_1, s => l8c7_0, cout => l8c8_0);
halfadder105: half_adder port map(x => l7c8_0, y => l7c8_1, s => l8c8_1, cout => l8c9_0);
halfadder106: half_adder port map(x => l7c9_0, y => l7c9_1, s => l8c9_1, cout => l8c10_0);
halfadder107: half_adder port map(x => l7c10_0, y => l7c10_1, s => l8c10_1, cout => l8c11_0);
halfadder108: half_adder port map(x => l7c11_0, y => l7c11_1, s => l8c11_1, cout => l8c12_0);
halfadder109: half_adder port map(x => l7c12_0, y => l7c12_1, s => l8c12_1, cout => l8c13_0);
halfadder110: half_adder port map(x => l7c13_0, y => l7c13_1, s => l8c13_1, cout => l8c14_0);
halfadder111: half_adder port map(x => l7c14_0, y => l7c14_1, s => l8c14_1, cout => l8c15_0);
halfadder112: half_adder port map(x => l7c15_0, y => l7c15_1, s => l8c15_1, cout => l8c16_0);
halfadder113: half_adder port map(x => l7c16_0, y => l7c16_1, s => l8c16_1, cout => l8c17_0);
halfadder114: half_adder port map(x => l7c17_0, y => l7c17_1, s => l8c17_1, cout => l8c18_0);
halfadder115: half_adder port map(x => l7c18_0, y => l7c18_1, s => l8c18_1, cout => l8c19_0);
halfadder116: half_adder port map(x => l7c19_0, y => l7c19_1, s => l8c19_1, cout => l8c20_0);
halfadder117: half_adder port map(x => l7c20_0, y => l7c20_1, s => l8c20_1, cout => l8c21_0);
halfadder118: half_adder port map(x => l7c21_0, y => l7c21_1, s => l8c21_1, cout => l8c22_0);
halfadder119: half_adder port map(x => l7c30_0, y => l7c30_1, s => l8c30_1, cout => l8c31_0);
halfadder120: half_adder port map(x => l7c31_0, y => l7c31_1, s => l8c31_1, cout => l8c32_0);
halfadder121: half_adder port map(x => l7c32_0, y => l7c32_1, s => l8c32_1, cout => l8c33_0);
halfadder122: half_adder port map(x => l7c33_0, y => l7c33_1, s => l8c33_1, cout => l8c34_0);
halfadder123: half_adder port map(x => l7c34_0, y => l7c34_1, s => l8c34_1, cout => l8c35_0);
halfadder124: half_adder port map(x => l7c35_0, y => l7c35_1, s => l8c35_1, cout => l8c36_0);
halfadder125: half_adder port map(x => l7c36_0, y => l7c36_1, s => l8c36_1, cout => l8c37_0);
halfadder126: half_adder port map(x => l7c37_0, y => l7c37_1, s => l8c37_1, cout => l8c38_0);
halfadder127: half_adder port map(x => l7c38_0, y => l7c38_1, s => l8c38_1, cout => l8c39_0);
halfadder128: half_adder port map(x => l7c39_0, y => l7c39_1, s => l8c39_1, cout => l8c40_0);
halfadder129: half_adder port map(x => l7c40_0, y => l7c40_1, s => l8c40_1, cout => l8c41_0);
halfadder130: half_adder port map(x => l7c41_0, y => l7c41_1, s => l8c41_1, cout => l8c42_0);
halfadder131: half_adder port map(x => l7c42_0, y => l7c42_1, s => l8c42_1, cout => l8c43_0);
halfadder132: half_adder port map(x => l7c43_0, y => l7c43_1, s => l8c43_1, cout => l8c44_0);
halfadder133: half_adder port map(x => l7c44_0, y => l7c44_1, s => l8c44_1, cout => l8c45_0);
halfadder134: half_adder port map(x => l7c45_0, y => l7c45_1, s => l8c45_1, cout => l8c46_0);
halfadder135: half_adder port map(x => l7c46_0, y => l7c46_1, s => l8c46_1, cout => l8c47_0);
halfadder136: half_adder port map(x => l7c47_0, y => l7c47_1, s => l8c47_1, cout => l8c48_0);

fulladder0: full_adder port map(x => l1c2_0, y => l1c2_1, cin => l1c2_2, s => l2c2_1, cout => l2c3_0);
fulladder1: full_adder port map(x => l1c3_0, y => l1c3_1, cin => l1c3_2, s => l2c3_1, cout => l2c4_0);
fulladder2: full_adder port map(x => l1c4_0, y => l1c4_1, cin => l1c4_2, s => l2c4_1, cout => l2c5_0);
fulladder3: full_adder port map(x => l1c5_0, y => l1c5_1, cin => l1c5_2, s => l2c5_2, cout => l2c6_0);
fulladder4: full_adder port map(x => l1c5_3, y => l1c5_4, cin => l1c5_5, s => l2c5_3, cout => l2c6_1);
fulladder5: full_adder port map(x => l1c6_0, y => l1c6_1, cin => l1c6_2, s => l2c6_2, cout => l2c7_0);
fulladder6: full_adder port map(x => l1c6_3, y => l1c6_4, cin => l1c6_5, s => l2c6_3, cout => l2c7_1);
fulladder7: full_adder port map(x => l1c7_0, y => l1c7_1, cin => l1c7_2, s => l2c7_2, cout => l2c8_0);
fulladder8: full_adder port map(x => l1c7_3, y => l1c7_4, cin => l1c7_5, s => l2c7_3, cout => l2c8_1);
fulladder9: full_adder port map(x => l1c8_0, y => l1c8_1, cin => l1c8_2, s => l2c8_3, cout => l2c9_0);
fulladder10: full_adder port map(x => l1c8_3, y => l1c8_4, cin => l1c8_5, s => l2c8_4, cout => l2c9_1);
fulladder11: full_adder port map(x => l1c8_6, y => l1c8_7, cin => l1c8_8, s => l2c8_5, cout => l2c9_2);
fulladder12: full_adder port map(x => l1c9_0, y => l1c9_1, cin => l1c9_2, s => l2c9_3, cout => l2c10_0);
fulladder13: full_adder port map(x => l1c9_3, y => l1c9_4, cin => l1c9_5, s => l2c9_4, cout => l2c10_1);
fulladder14: full_adder port map(x => l1c9_6, y => l1c9_7, cin => l1c9_8, s => l2c9_5, cout => l2c10_2);
fulladder15: full_adder port map(x => l1c10_0, y => l1c10_1, cin => l1c10_2, s => l2c10_3, cout => l2c11_0);
fulladder16: full_adder port map(x => l1c10_3, y => l1c10_4, cin => l1c10_5, s => l2c10_4, cout => l2c11_1);
fulladder17: full_adder port map(x => l1c10_6, y => l1c10_7, cin => l1c10_8, s => l2c10_5, cout => l2c11_2);
fulladder18: full_adder port map(x => l1c11_0, y => l1c11_1, cin => l1c11_2, s => l2c11_4, cout => l2c12_0);
fulladder19: full_adder port map(x => l1c11_3, y => l1c11_4, cin => l1c11_5, s => l2c11_5, cout => l2c12_1);
fulladder20: full_adder port map(x => l1c11_6, y => l1c11_7, cin => l1c11_8, s => l2c11_6, cout => l2c12_2);
fulladder21: full_adder port map(x => l1c11_9, y => l1c11_10, cin => l1c11_11, s => l2c11_7, cout => l2c12_3);
fulladder22: full_adder port map(x => l1c12_0, y => l1c12_1, cin => l1c12_2, s => l2c12_4, cout => l2c13_0);
fulladder23: full_adder port map(x => l1c12_3, y => l1c12_4, cin => l1c12_5, s => l2c12_5, cout => l2c13_1);
fulladder24: full_adder port map(x => l1c12_6, y => l1c12_7, cin => l1c12_8, s => l2c12_6, cout => l2c13_2);
fulladder25: full_adder port map(x => l1c12_9, y => l1c12_10, cin => l1c12_11, s => l2c12_7, cout => l2c13_3);
fulladder26: full_adder port map(x => l1c13_0, y => l1c13_1, cin => l1c13_2, s => l2c13_4, cout => l2c14_0);
fulladder27: full_adder port map(x => l1c13_3, y => l1c13_4, cin => l1c13_5, s => l2c13_5, cout => l2c14_1);
fulladder28: full_adder port map(x => l1c13_6, y => l1c13_7, cin => l1c13_8, s => l2c13_6, cout => l2c14_2);
fulladder29: full_adder port map(x => l1c13_9, y => l1c13_10, cin => l1c13_11, s => l2c13_7, cout => l2c14_3);
fulladder30: full_adder port map(x => l1c14_0, y => l1c14_1, cin => l1c14_2, s => l2c14_5, cout => l2c15_0);
fulladder31: full_adder port map(x => l1c14_3, y => l1c14_4, cin => l1c14_5, s => l2c14_6, cout => l2c15_1);
fulladder32: full_adder port map(x => l1c14_6, y => l1c14_7, cin => l1c14_8, s => l2c14_7, cout => l2c15_2);
fulladder33: full_adder port map(x => l1c14_9, y => l1c14_10, cin => l1c14_11, s => l2c14_8, cout => l2c15_3);
fulladder34: full_adder port map(x => l1c14_12, y => l1c14_13, cin => l1c14_14, s => l2c14_9, cout => l2c15_4);
fulladder35: full_adder port map(x => l1c15_0, y => l1c15_1, cin => l1c15_2, s => l2c15_5, cout => l2c16_0);
fulladder36: full_adder port map(x => l1c15_3, y => l1c15_4, cin => l1c15_5, s => l2c15_6, cout => l2c16_1);
fulladder37: full_adder port map(x => l1c15_6, y => l1c15_7, cin => l1c15_8, s => l2c15_7, cout => l2c16_2);
fulladder38: full_adder port map(x => l1c15_9, y => l1c15_10, cin => l1c15_11, s => l2c15_8, cout => l2c16_3);
fulladder39: full_adder port map(x => l1c15_12, y => l1c15_13, cin => l1c15_14, s => l2c15_9, cout => l2c16_4);
fulladder40: full_adder port map(x => l1c16_0, y => l1c16_1, cin => l1c16_2, s => l2c16_5, cout => l2c17_0);
fulladder41: full_adder port map(x => l1c16_3, y => l1c16_4, cin => l1c16_5, s => l2c16_6, cout => l2c17_1);
fulladder42: full_adder port map(x => l1c16_6, y => l1c16_7, cin => l1c16_8, s => l2c16_7, cout => l2c17_2);
fulladder43: full_adder port map(x => l1c16_9, y => l1c16_10, cin => l1c16_11, s => l2c16_8, cout => l2c17_3);
fulladder44: full_adder port map(x => l1c16_12, y => l1c16_13, cin => l1c16_14, s => l2c16_9, cout => l2c17_4);
fulladder45: full_adder port map(x => l1c17_0, y => l1c17_1, cin => l1c17_2, s => l2c17_6, cout => l2c18_0);
fulladder46: full_adder port map(x => l1c17_3, y => l1c17_4, cin => l1c17_5, s => l2c17_7, cout => l2c18_1);
fulladder47: full_adder port map(x => l1c17_6, y => l1c17_7, cin => l1c17_8, s => l2c17_8, cout => l2c18_2);
fulladder48: full_adder port map(x => l1c17_9, y => l1c17_10, cin => l1c17_11, s => l2c17_9, cout => l2c18_3);
fulladder49: full_adder port map(x => l1c17_12, y => l1c17_13, cin => l1c17_14, s => l2c17_10, cout => l2c18_4);
fulladder50: full_adder port map(x => l1c17_15, y => l1c17_16, cin => l1c17_17, s => l2c17_11, cout => l2c18_5);
fulladder51: full_adder port map(x => l1c18_0, y => l1c18_1, cin => l1c18_2, s => l2c18_6, cout => l2c19_0);
fulladder52: full_adder port map(x => l1c18_3, y => l1c18_4, cin => l1c18_5, s => l2c18_7, cout => l2c19_1);
fulladder53: full_adder port map(x => l1c18_6, y => l1c18_7, cin => l1c18_8, s => l2c18_8, cout => l2c19_2);
fulladder54: full_adder port map(x => l1c18_9, y => l1c18_10, cin => l1c18_11, s => l2c18_9, cout => l2c19_3);
fulladder55: full_adder port map(x => l1c18_12, y => l1c18_13, cin => l1c18_14, s => l2c18_10, cout => l2c19_4);
fulladder56: full_adder port map(x => l1c18_15, y => l1c18_16, cin => l1c18_17, s => l2c18_11, cout => l2c19_5);
fulladder57: full_adder port map(x => l1c19_0, y => l1c19_1, cin => l1c19_2, s => l2c19_6, cout => l2c20_0);
fulladder58: full_adder port map(x => l1c19_3, y => l1c19_4, cin => l1c19_5, s => l2c19_7, cout => l2c20_1);
fulladder59: full_adder port map(x => l1c19_6, y => l1c19_7, cin => l1c19_8, s => l2c19_8, cout => l2c20_2);
fulladder60: full_adder port map(x => l1c19_9, y => l1c19_10, cin => l1c19_11, s => l2c19_9, cout => l2c20_3);
fulladder61: full_adder port map(x => l1c19_12, y => l1c19_13, cin => l1c19_14, s => l2c19_10, cout => l2c20_4);
fulladder62: full_adder port map(x => l1c19_15, y => l1c19_16, cin => l1c19_17, s => l2c19_11, cout => l2c20_5);
fulladder63: full_adder port map(x => l1c20_0, y => l1c20_1, cin => l1c20_2, s => l2c20_7, cout => l2c21_0);
fulladder64: full_adder port map(x => l1c20_3, y => l1c20_4, cin => l1c20_5, s => l2c20_8, cout => l2c21_1);
fulladder65: full_adder port map(x => l1c20_6, y => l1c20_7, cin => l1c20_8, s => l2c20_9, cout => l2c21_2);
fulladder66: full_adder port map(x => l1c20_9, y => l1c20_10, cin => l1c20_11, s => l2c20_10, cout => l2c21_3);
fulladder67: full_adder port map(x => l1c20_12, y => l1c20_13, cin => l1c20_14, s => l2c20_11, cout => l2c21_4);
fulladder68: full_adder port map(x => l1c20_15, y => l1c20_16, cin => l1c20_17, s => l2c20_12, cout => l2c21_5);
fulladder69: full_adder port map(x => l1c20_18, y => l1c20_19, cin => l1c20_20, s => l2c20_13, cout => l2c21_6);
fulladder70: full_adder port map(x => l1c21_0, y => l1c21_1, cin => l1c21_2, s => l2c21_7, cout => l2c22_0);
fulladder71: full_adder port map(x => l1c21_3, y => l1c21_4, cin => l1c21_5, s => l2c21_8, cout => l2c22_1);
fulladder72: full_adder port map(x => l1c21_6, y => l1c21_7, cin => l1c21_8, s => l2c21_9, cout => l2c22_2);
fulladder73: full_adder port map(x => l1c21_9, y => l1c21_10, cin => l1c21_11, s => l2c21_10, cout => l2c22_3);
fulladder74: full_adder port map(x => l1c21_12, y => l1c21_13, cin => l1c21_14, s => l2c21_11, cout => l2c22_4);
fulladder75: full_adder port map(x => l1c21_15, y => l1c21_16, cin => l1c21_17, s => l2c21_12, cout => l2c22_5);
fulladder76: full_adder port map(x => l1c21_18, y => l1c21_19, cin => l1c21_20, s => l2c21_13, cout => l2c22_6);
fulladder77: full_adder port map(x => l1c22_0, y => l1c22_1, cin => l1c22_2, s => l2c22_7, cout => l2c23_0);
fulladder78: full_adder port map(x => l1c22_3, y => l1c22_4, cin => l1c22_5, s => l2c22_8, cout => l2c23_1);
fulladder79: full_adder port map(x => l1c22_6, y => l1c22_7, cin => l1c22_8, s => l2c22_9, cout => l2c23_2);
fulladder80: full_adder port map(x => l1c22_9, y => l1c22_10, cin => l1c22_11, s => l2c22_10, cout => l2c23_3);
fulladder81: full_adder port map(x => l1c22_12, y => l1c22_13, cin => l1c22_14, s => l2c22_11, cout => l2c23_4);
fulladder82: full_adder port map(x => l1c22_15, y => l1c22_16, cin => l1c22_17, s => l2c22_12, cout => l2c23_5);
fulladder83: full_adder port map(x => l1c22_18, y => l1c22_19, cin => l1c22_20, s => l2c22_13, cout => l2c23_6);
fulladder84: full_adder port map(x => l1c23_0, y => l1c23_1, cin => l1c23_2, s => l2c23_8, cout => l2c24_0);
fulladder85: full_adder port map(x => l1c23_3, y => l1c23_4, cin => l1c23_5, s => l2c23_9, cout => l2c24_1);
fulladder86: full_adder port map(x => l1c23_6, y => l1c23_7, cin => l1c23_8, s => l2c23_10, cout => l2c24_2);
fulladder87: full_adder port map(x => l1c23_9, y => l1c23_10, cin => l1c23_11, s => l2c23_11, cout => l2c24_3);
fulladder88: full_adder port map(x => l1c23_12, y => l1c23_13, cin => l1c23_14, s => l2c23_12, cout => l2c24_4);
fulladder89: full_adder port map(x => l1c23_15, y => l1c23_16, cin => l1c23_17, s => l2c23_13, cout => l2c24_5);
fulladder90: full_adder port map(x => l1c23_18, y => l1c23_19, cin => l1c23_20, s => l2c23_14, cout => l2c24_6);
fulladder91: full_adder port map(x => l1c23_21, y => l1c23_22, cin => l1c23_23, s => l2c23_15, cout => l2c24_7);
fulladder92: full_adder port map(x => l1c24_0, y => l1c24_1, cin => l1c24_2, s => l2c24_8, cout => l2c25_0);
fulladder93: full_adder port map(x => l1c24_3, y => l1c24_4, cin => l1c24_5, s => l2c24_9, cout => l2c25_1);
fulladder94: full_adder port map(x => l1c24_6, y => l1c24_7, cin => l1c24_8, s => l2c24_10, cout => l2c25_2);
fulladder95: full_adder port map(x => l1c24_9, y => l1c24_10, cin => l1c24_11, s => l2c24_11, cout => l2c25_3);
fulladder96: full_adder port map(x => l1c24_12, y => l1c24_13, cin => l1c24_14, s => l2c24_12, cout => l2c25_4);
fulladder97: full_adder port map(x => l1c24_15, y => l1c24_16, cin => l1c24_17, s => l2c24_13, cout => l2c25_5);
fulladder98: full_adder port map(x => l1c24_18, y => l1c24_19, cin => l1c24_20, s => l2c24_14, cout => l2c25_6);
fulladder99: full_adder port map(x => l1c25_0, y => l1c25_1, cin => l1c25_2, s => l2c25_8, cout => l2c26_0);
fulladder100: full_adder port map(x => l1c25_3, y => l1c25_4, cin => l1c25_5, s => l2c25_9, cout => l2c26_1);
fulladder101: full_adder port map(x => l1c25_6, y => l1c25_7, cin => l1c25_8, s => l2c25_10, cout => l2c26_2);
fulladder102: full_adder port map(x => l1c25_9, y => l1c25_10, cin => l1c25_11, s => l2c25_11, cout => l2c26_3);
fulladder103: full_adder port map(x => l1c25_12, y => l1c25_13, cin => l1c25_14, s => l2c25_12, cout => l2c26_4);
fulladder104: full_adder port map(x => l1c25_15, y => l1c25_16, cin => l1c25_17, s => l2c25_13, cout => l2c26_5);
fulladder105: full_adder port map(x => l1c25_18, y => l1c25_19, cin => l1c25_20, s => l2c25_14, cout => l2c26_6);
fulladder106: full_adder port map(x => l1c26_0, y => l1c26_1, cin => l1c26_2, s => l2c26_7, cout => l2c27_0);
fulladder107: full_adder port map(x => l1c26_3, y => l1c26_4, cin => l1c26_5, s => l2c26_8, cout => l2c27_1);
fulladder108: full_adder port map(x => l1c26_6, y => l1c26_7, cin => l1c26_8, s => l2c26_9, cout => l2c27_2);
fulladder109: full_adder port map(x => l1c26_9, y => l1c26_10, cin => l1c26_11, s => l2c26_10, cout => l2c27_3);
fulladder110: full_adder port map(x => l1c26_12, y => l1c26_13, cin => l1c26_14, s => l2c26_11, cout => l2c27_4);
fulladder111: full_adder port map(x => l1c26_15, y => l1c26_16, cin => l1c26_17, s => l2c26_12, cout => l2c27_5);
fulladder112: full_adder port map(x => l1c26_18, y => l1c26_19, cin => l1c26_20, s => l2c26_13, cout => l2c27_6);
fulladder113: full_adder port map(x => l1c27_0, y => l1c27_1, cin => l1c27_2, s => l2c27_7, cout => l2c28_0);
fulladder114: full_adder port map(x => l1c27_3, y => l1c27_4, cin => l1c27_5, s => l2c27_8, cout => l2c28_1);
fulladder115: full_adder port map(x => l1c27_6, y => l1c27_7, cin => l1c27_8, s => l2c27_9, cout => l2c28_2);
fulladder116: full_adder port map(x => l1c27_9, y => l1c27_10, cin => l1c27_11, s => l2c27_10, cout => l2c28_3);
fulladder117: full_adder port map(x => l1c27_12, y => l1c27_13, cin => l1c27_14, s => l2c27_11, cout => l2c28_4);
fulladder118: full_adder port map(x => l1c27_15, y => l1c27_16, cin => l1c27_17, s => l2c27_12, cout => l2c28_5);
fulladder119: full_adder port map(x => l1c28_0, y => l1c28_1, cin => l1c28_2, s => l2c28_7, cout => l2c29_0);
fulladder120: full_adder port map(x => l1c28_3, y => l1c28_4, cin => l1c28_5, s => l2c28_8, cout => l2c29_1);
fulladder121: full_adder port map(x => l1c28_6, y => l1c28_7, cin => l1c28_8, s => l2c28_9, cout => l2c29_2);
fulladder122: full_adder port map(x => l1c28_9, y => l1c28_10, cin => l1c28_11, s => l2c28_10, cout => l2c29_3);
fulladder123: full_adder port map(x => l1c28_12, y => l1c28_13, cin => l1c28_14, s => l2c28_11, cout => l2c29_4);
fulladder124: full_adder port map(x => l1c28_15, y => l1c28_16, cin => l1c28_17, s => l2c28_12, cout => l2c29_5);
fulladder125: full_adder port map(x => l1c29_0, y => l1c29_1, cin => l1c29_2, s => l2c29_6, cout => l2c30_0);
fulladder126: full_adder port map(x => l1c29_3, y => l1c29_4, cin => l1c29_5, s => l2c29_7, cout => l2c30_1);
fulladder127: full_adder port map(x => l1c29_6, y => l1c29_7, cin => l1c29_8, s => l2c29_8, cout => l2c30_2);
fulladder128: full_adder port map(x => l1c29_9, y => l1c29_10, cin => l1c29_11, s => l2c29_9, cout => l2c30_3);
fulladder129: full_adder port map(x => l1c29_12, y => l1c29_13, cin => l1c29_14, s => l2c29_10, cout => l2c30_4);
fulladder130: full_adder port map(x => l1c29_15, y => l1c29_16, cin => l1c29_17, s => l2c29_11, cout => l2c30_5);
fulladder131: full_adder port map(x => l1c30_0, y => l1c30_1, cin => l1c30_2, s => l2c30_6, cout => l2c31_0);
fulladder132: full_adder port map(x => l1c30_3, y => l1c30_4, cin => l1c30_5, s => l2c30_7, cout => l2c31_1);
fulladder133: full_adder port map(x => l1c30_6, y => l1c30_7, cin => l1c30_8, s => l2c30_8, cout => l2c31_2);
fulladder134: full_adder port map(x => l1c30_9, y => l1c30_10, cin => l1c30_11, s => l2c30_9, cout => l2c31_3);
fulladder135: full_adder port map(x => l1c30_12, y => l1c30_13, cin => l1c30_14, s => l2c30_10, cout => l2c31_4);
fulladder136: full_adder port map(x => l1c31_0, y => l1c31_1, cin => l1c31_2, s => l2c31_6, cout => l2c32_0);
fulladder137: full_adder port map(x => l1c31_3, y => l1c31_4, cin => l1c31_5, s => l2c31_7, cout => l2c32_1);
fulladder138: full_adder port map(x => l1c31_6, y => l1c31_7, cin => l1c31_8, s => l2c31_8, cout => l2c32_2);
fulladder139: full_adder port map(x => l1c31_9, y => l1c31_10, cin => l1c31_11, s => l2c31_9, cout => l2c32_3);
fulladder140: full_adder port map(x => l1c31_12, y => l1c31_13, cin => l1c31_14, s => l2c31_10, cout => l2c32_4);
fulladder141: full_adder port map(x => l1c32_0, y => l1c32_1, cin => l1c32_2, s => l2c32_5, cout => l2c33_0);
fulladder142: full_adder port map(x => l1c32_3, y => l1c32_4, cin => l1c32_5, s => l2c32_6, cout => l2c33_1);
fulladder143: full_adder port map(x => l1c32_6, y => l1c32_7, cin => l1c32_8, s => l2c32_7, cout => l2c33_2);
fulladder144: full_adder port map(x => l1c32_9, y => l1c32_10, cin => l1c32_11, s => l2c32_8, cout => l2c33_3);
fulladder145: full_adder port map(x => l1c32_12, y => l1c32_13, cin => l1c32_14, s => l2c32_9, cout => l2c33_4);
fulladder146: full_adder port map(x => l1c33_0, y => l1c33_1, cin => l1c33_2, s => l2c33_5, cout => l2c34_0);
fulladder147: full_adder port map(x => l1c33_3, y => l1c33_4, cin => l1c33_5, s => l2c33_6, cout => l2c34_1);
fulladder148: full_adder port map(x => l1c33_6, y => l1c33_7, cin => l1c33_8, s => l2c33_7, cout => l2c34_2);
fulladder149: full_adder port map(x => l1c33_9, y => l1c33_10, cin => l1c33_11, s => l2c33_8, cout => l2c34_3);
fulladder150: full_adder port map(x => l1c34_0, y => l1c34_1, cin => l1c34_2, s => l2c34_5, cout => l2c35_0);
fulladder151: full_adder port map(x => l1c34_3, y => l1c34_4, cin => l1c34_5, s => l2c34_6, cout => l2c35_1);
fulladder152: full_adder port map(x => l1c34_6, y => l1c34_7, cin => l1c34_8, s => l2c34_7, cout => l2c35_2);
fulladder153: full_adder port map(x => l1c34_9, y => l1c34_10, cin => l1c34_11, s => l2c34_8, cout => l2c35_3);
fulladder154: full_adder port map(x => l1c35_0, y => l1c35_1, cin => l1c35_2, s => l2c35_4, cout => l2c36_0);
fulladder155: full_adder port map(x => l1c35_3, y => l1c35_4, cin => l1c35_5, s => l2c35_5, cout => l2c36_1);
fulladder156: full_adder port map(x => l1c35_6, y => l1c35_7, cin => l1c35_8, s => l2c35_6, cout => l2c36_2);
fulladder157: full_adder port map(x => l1c35_9, y => l1c35_10, cin => l1c35_11, s => l2c35_7, cout => l2c36_3);
fulladder158: full_adder port map(x => l1c36_0, y => l1c36_1, cin => l1c36_2, s => l2c36_4, cout => l2c37_0);
fulladder159: full_adder port map(x => l1c36_3, y => l1c36_4, cin => l1c36_5, s => l2c36_5, cout => l2c37_1);
fulladder160: full_adder port map(x => l1c36_6, y => l1c36_7, cin => l1c36_8, s => l2c36_6, cout => l2c37_2);
fulladder161: full_adder port map(x => l1c37_0, y => l1c37_1, cin => l1c37_2, s => l2c37_4, cout => l2c38_0);
fulladder162: full_adder port map(x => l1c37_3, y => l1c37_4, cin => l1c37_5, s => l2c37_5, cout => l2c38_1);
fulladder163: full_adder port map(x => l1c37_6, y => l1c37_7, cin => l1c37_8, s => l2c37_6, cout => l2c38_2);
fulladder164: full_adder port map(x => l1c38_0, y => l1c38_1, cin => l1c38_2, s => l2c38_3, cout => l2c39_0);
fulladder165: full_adder port map(x => l1c38_3, y => l1c38_4, cin => l1c38_5, s => l2c38_4, cout => l2c39_1);
fulladder166: full_adder port map(x => l1c38_6, y => l1c38_7, cin => l1c38_8, s => l2c38_5, cout => l2c39_2);
fulladder167: full_adder port map(x => l1c39_0, y => l1c39_1, cin => l1c39_2, s => l2c39_3, cout => l2c40_0);
fulladder168: full_adder port map(x => l1c39_3, y => l1c39_4, cin => l1c39_5, s => l2c39_4, cout => l2c40_1);
fulladder169: full_adder port map(x => l1c40_0, y => l1c40_1, cin => l1c40_2, s => l2c40_3, cout => l2c41_0);
fulladder170: full_adder port map(x => l1c40_3, y => l1c40_4, cin => l1c40_5, s => l2c40_4, cout => l2c41_1);
fulladder171: full_adder port map(x => l1c41_0, y => l1c41_1, cin => l1c41_2, s => l2c41_2, cout => l2c42_0);
fulladder172: full_adder port map(x => l1c41_3, y => l1c41_4, cin => l1c41_5, s => l2c41_3, cout => l2c42_1);
fulladder173: full_adder port map(x => l1c42_0, y => l1c42_1, cin => l1c42_2, s => l2c42_2, cout => l2c43_0);
fulladder174: full_adder port map(x => l1c43_0, y => l1c43_1, cin => l1c43_2, s => l2c43_2, cout => l2c44_0);
fulladder175: full_adder port map(x => l1c44_0, y => l1c44_1, cin => l1c44_2, s => l2c44_1, cout => l2c45_0);
fulladder176: full_adder port map(x => l2c3_0, y => l2c3_1, cin => l1c3_3, s => l3c3_1, cout => l3c4_0);
fulladder177: full_adder port map(x => l2c4_0, y => l2c4_1, cin => l2c4_2, s => l3c4_1, cout => l3c5_0);
fulladder178: full_adder port map(x => l2c5_0, y => l2c5_1, cin => l2c5_2, s => l3c5_1, cout => l3c6_0);
fulladder179: full_adder port map(x => l2c6_0, y => l2c6_1, cin => l2c6_2, s => l3c6_1, cout => l3c7_0);
fulladder180: full_adder port map(x => l2c7_0, y => l2c7_1, cin => l2c7_2, s => l3c7_2, cout => l3c8_0);
fulladder181: full_adder port map(x => l2c8_0, y => l2c8_1, cin => l2c8_2, s => l3c8_2, cout => l3c9_0);
fulladder182: full_adder port map(x => l2c8_3, y => l2c8_4, cin => l2c8_5, s => l3c8_3, cout => l3c9_1);
fulladder183: full_adder port map(x => l2c9_0, y => l2c9_1, cin => l2c9_2, s => l3c9_2, cout => l3c10_0);
fulladder184: full_adder port map(x => l2c9_3, y => l2c9_4, cin => l2c9_5, s => l3c9_3, cout => l3c10_1);
fulladder185: full_adder port map(x => l2c10_0, y => l2c10_1, cin => l2c10_2, s => l3c10_2, cout => l3c11_0);
fulladder186: full_adder port map(x => l2c10_3, y => l2c10_4, cin => l2c10_5, s => l3c10_3, cout => l3c11_1);
fulladder187: full_adder port map(x => l2c11_0, y => l2c11_1, cin => l2c11_2, s => l3c11_2, cout => l3c12_0);
fulladder188: full_adder port map(x => l2c11_3, y => l2c11_4, cin => l2c11_5, s => l3c11_3, cout => l3c12_1);
fulladder189: full_adder port map(x => l2c12_0, y => l2c12_1, cin => l2c12_2, s => l3c12_3, cout => l3c13_0);
fulladder190: full_adder port map(x => l2c12_3, y => l2c12_4, cin => l2c12_5, s => l3c12_4, cout => l3c13_1);
fulladder191: full_adder port map(x => l2c12_6, y => l2c12_7, cin => l1c12_12, s => l3c12_5, cout => l3c13_2);
fulladder192: full_adder port map(x => l2c13_0, y => l2c13_1, cin => l2c13_2, s => l3c13_3, cout => l3c14_0);
fulladder193: full_adder port map(x => l2c13_3, y => l2c13_4, cin => l2c13_5, s => l3c13_4, cout => l3c14_1);
fulladder194: full_adder port map(x => l2c13_6, y => l2c13_7, cin => l2c13_8, s => l3c13_5, cout => l3c14_2);
fulladder195: full_adder port map(x => l2c14_0, y => l2c14_1, cin => l2c14_2, s => l3c14_3, cout => l3c15_0);
fulladder196: full_adder port map(x => l2c14_3, y => l2c14_4, cin => l2c14_5, s => l3c14_4, cout => l3c15_1);
fulladder197: full_adder port map(x => l2c14_6, y => l2c14_7, cin => l2c14_8, s => l3c14_5, cout => l3c15_2);
fulladder198: full_adder port map(x => l2c15_0, y => l2c15_1, cin => l2c15_2, s => l3c15_3, cout => l3c16_0);
fulladder199: full_adder port map(x => l2c15_3, y => l2c15_4, cin => l2c15_5, s => l3c15_4, cout => l3c16_1);
fulladder200: full_adder port map(x => l2c15_6, y => l2c15_7, cin => l2c15_8, s => l3c15_5, cout => l3c16_2);
fulladder201: full_adder port map(x => l2c16_0, y => l2c16_1, cin => l2c16_2, s => l3c16_4, cout => l3c17_0);
fulladder202: full_adder port map(x => l2c16_3, y => l2c16_4, cin => l2c16_5, s => l3c16_5, cout => l3c17_1);
fulladder203: full_adder port map(x => l2c16_6, y => l2c16_7, cin => l2c16_8, s => l3c16_6, cout => l3c17_2);
fulladder204: full_adder port map(x => l2c17_0, y => l2c17_1, cin => l2c17_2, s => l3c17_4, cout => l3c18_0);
fulladder205: full_adder port map(x => l2c17_3, y => l2c17_4, cin => l2c17_5, s => l3c17_5, cout => l3c18_1);
fulladder206: full_adder port map(x => l2c17_6, y => l2c17_7, cin => l2c17_8, s => l3c17_6, cout => l3c18_2);
fulladder207: full_adder port map(x => l2c17_9, y => l2c17_10, cin => l2c17_11, s => l3c17_7, cout => l3c18_3);
fulladder208: full_adder port map(x => l2c18_0, y => l2c18_1, cin => l2c18_2, s => l3c18_4, cout => l3c19_0);
fulladder209: full_adder port map(x => l2c18_3, y => l2c18_4, cin => l2c18_5, s => l3c18_5, cout => l3c19_1);
fulladder210: full_adder port map(x => l2c18_6, y => l2c18_7, cin => l2c18_8, s => l3c18_6, cout => l3c19_2);
fulladder211: full_adder port map(x => l2c18_9, y => l2c18_10, cin => l2c18_11, s => l3c18_7, cout => l3c19_3);
fulladder212: full_adder port map(x => l2c19_0, y => l2c19_1, cin => l2c19_2, s => l3c19_4, cout => l3c20_0);
fulladder213: full_adder port map(x => l2c19_3, y => l2c19_4, cin => l2c19_5, s => l3c19_5, cout => l3c20_1);
fulladder214: full_adder port map(x => l2c19_6, y => l2c19_7, cin => l2c19_8, s => l3c19_6, cout => l3c20_2);
fulladder215: full_adder port map(x => l2c19_9, y => l2c19_10, cin => l2c19_11, s => l3c19_7, cout => l3c20_3);
fulladder216: full_adder port map(x => l2c20_0, y => l2c20_1, cin => l2c20_2, s => l3c20_4, cout => l3c21_0);
fulladder217: full_adder port map(x => l2c20_3, y => l2c20_4, cin => l2c20_5, s => l3c20_5, cout => l3c21_1);
fulladder218: full_adder port map(x => l2c20_6, y => l2c20_7, cin => l2c20_8, s => l3c20_6, cout => l3c21_2);
fulladder219: full_adder port map(x => l2c20_9, y => l2c20_10, cin => l2c20_11, s => l3c20_7, cout => l3c21_3);
fulladder220: full_adder port map(x => l2c21_0, y => l2c21_1, cin => l2c21_2, s => l3c21_5, cout => l3c22_0);
fulladder221: full_adder port map(x => l2c21_3, y => l2c21_4, cin => l2c21_5, s => l3c21_6, cout => l3c22_1);
fulladder222: full_adder port map(x => l2c21_6, y => l2c21_7, cin => l2c21_8, s => l3c21_7, cout => l3c22_2);
fulladder223: full_adder port map(x => l2c21_9, y => l2c21_10, cin => l2c21_11, s => l3c21_8, cout => l3c22_3);
fulladder224: full_adder port map(x => l2c21_12, y => l2c21_13, cin => l1c21_21, s => l3c21_9, cout => l3c22_4);
fulladder225: full_adder port map(x => l2c22_0, y => l2c22_1, cin => l2c22_2, s => l3c22_5, cout => l3c23_0);
fulladder226: full_adder port map(x => l2c22_3, y => l2c22_4, cin => l2c22_5, s => l3c22_6, cout => l3c23_1);
fulladder227: full_adder port map(x => l2c22_6, y => l2c22_7, cin => l2c22_8, s => l3c22_7, cout => l3c23_2);
fulladder228: full_adder port map(x => l2c22_9, y => l2c22_10, cin => l2c22_11, s => l3c22_8, cout => l3c23_3);
fulladder229: full_adder port map(x => l2c22_12, y => l2c22_13, cin => l2c22_14, s => l3c22_9, cout => l3c23_4);
fulladder230: full_adder port map(x => l2c23_0, y => l2c23_1, cin => l2c23_2, s => l3c23_5, cout => l3c24_0);
fulladder231: full_adder port map(x => l2c23_3, y => l2c23_4, cin => l2c23_5, s => l3c23_6, cout => l3c24_1);
fulladder232: full_adder port map(x => l2c23_6, y => l2c23_7, cin => l2c23_8, s => l3c23_7, cout => l3c24_2);
fulladder233: full_adder port map(x => l2c23_9, y => l2c23_10, cin => l2c23_11, s => l3c23_8, cout => l3c24_3);
fulladder234: full_adder port map(x => l2c23_12, y => l2c23_13, cin => l2c23_14, s => l3c23_9, cout => l3c24_4);
fulladder235: full_adder port map(x => l2c24_0, y => l2c24_1, cin => l2c24_2, s => l3c24_5, cout => l3c25_0);
fulladder236: full_adder port map(x => l2c24_3, y => l2c24_4, cin => l2c24_5, s => l3c24_6, cout => l3c25_1);
fulladder237: full_adder port map(x => l2c24_6, y => l2c24_7, cin => l2c24_8, s => l3c24_7, cout => l3c25_2);
fulladder238: full_adder port map(x => l2c24_9, y => l2c24_10, cin => l2c24_11, s => l3c24_8, cout => l3c25_3);
fulladder239: full_adder port map(x => l2c24_12, y => l2c24_13, cin => l2c24_14, s => l3c24_9, cout => l3c25_4);
fulladder240: full_adder port map(x => l2c25_0, y => l2c25_1, cin => l2c25_2, s => l3c25_5, cout => l3c26_0);
fulladder241: full_adder port map(x => l2c25_3, y => l2c25_4, cin => l2c25_5, s => l3c25_6, cout => l3c26_1);
fulladder242: full_adder port map(x => l2c25_6, y => l2c25_7, cin => l2c25_8, s => l3c25_7, cout => l3c26_2);
fulladder243: full_adder port map(x => l2c25_9, y => l2c25_10, cin => l2c25_11, s => l3c25_8, cout => l3c26_3);
fulladder244: full_adder port map(x => l2c25_12, y => l2c25_13, cin => l2c25_14, s => l3c25_9, cout => l3c26_4);
fulladder245: full_adder port map(x => l2c26_0, y => l2c26_1, cin => l2c26_2, s => l3c26_5, cout => l3c27_0);
fulladder246: full_adder port map(x => l2c26_3, y => l2c26_4, cin => l2c26_5, s => l3c26_6, cout => l3c27_1);
fulladder247: full_adder port map(x => l2c26_6, y => l2c26_7, cin => l2c26_8, s => l3c26_7, cout => l3c27_2);
fulladder248: full_adder port map(x => l2c26_9, y => l2c26_10, cin => l2c26_11, s => l3c26_8, cout => l3c27_3);
fulladder249: full_adder port map(x => l2c27_0, y => l2c27_1, cin => l2c27_2, s => l3c27_5, cout => l3c28_0);
fulladder250: full_adder port map(x => l2c27_3, y => l2c27_4, cin => l2c27_5, s => l3c27_6, cout => l3c28_1);
fulladder251: full_adder port map(x => l2c27_6, y => l2c27_7, cin => l2c27_8, s => l3c27_7, cout => l3c28_2);
fulladder252: full_adder port map(x => l2c27_9, y => l2c27_10, cin => l2c27_11, s => l3c27_8, cout => l3c28_3);
fulladder253: full_adder port map(x => l2c28_0, y => l2c28_1, cin => l2c28_2, s => l3c28_5, cout => l3c29_0);
fulladder254: full_adder port map(x => l2c28_3, y => l2c28_4, cin => l2c28_5, s => l3c28_6, cout => l3c29_1);
fulladder255: full_adder port map(x => l2c28_6, y => l2c28_7, cin => l2c28_8, s => l3c28_7, cout => l3c29_2);
fulladder256: full_adder port map(x => l2c28_9, y => l2c28_10, cin => l2c28_11, s => l3c28_8, cout => l3c29_3);
fulladder257: full_adder port map(x => l2c29_0, y => l2c29_1, cin => l2c29_2, s => l3c29_5, cout => l3c30_0);
fulladder258: full_adder port map(x => l2c29_3, y => l2c29_4, cin => l2c29_5, s => l3c29_6, cout => l3c30_1);
fulladder259: full_adder port map(x => l2c29_6, y => l2c29_7, cin => l2c29_8, s => l3c29_7, cout => l3c30_2);
fulladder260: full_adder port map(x => l2c29_9, y => l2c29_10, cin => l2c29_11, s => l3c29_8, cout => l3c30_3);
fulladder261: full_adder port map(x => l2c30_0, y => l2c30_1, cin => l2c30_2, s => l3c30_4, cout => l3c31_0);
fulladder262: full_adder port map(x => l2c30_3, y => l2c30_4, cin => l2c30_5, s => l3c30_5, cout => l3c31_1);
fulladder263: full_adder port map(x => l2c30_6, y => l2c30_7, cin => l2c30_8, s => l3c30_6, cout => l3c31_2);
fulladder264: full_adder port map(x => l2c30_9, y => l2c30_10, cin => l2c30_11, s => l3c30_7, cout => l3c31_3);
fulladder265: full_adder port map(x => l2c31_0, y => l2c31_1, cin => l2c31_2, s => l3c31_4, cout => l3c32_0);
fulladder266: full_adder port map(x => l2c31_3, y => l2c31_4, cin => l2c31_5, s => l3c31_5, cout => l3c32_1);
fulladder267: full_adder port map(x => l2c31_6, y => l2c31_7, cin => l2c31_8, s => l3c31_6, cout => l3c32_2);
fulladder268: full_adder port map(x => l2c31_9, y => l2c31_10, cin => l1c31_15, s => l3c31_7, cout => l3c32_3);
fulladder269: full_adder port map(x => l2c32_0, y => l2c32_1, cin => l2c32_2, s => l3c32_4, cout => l3c33_0);
fulladder270: full_adder port map(x => l2c32_3, y => l2c32_4, cin => l2c32_5, s => l3c32_5, cout => l3c33_1);
fulladder271: full_adder port map(x => l2c32_6, y => l2c32_7, cin => l2c32_8, s => l3c32_6, cout => l3c33_2);
fulladder272: full_adder port map(x => l2c33_0, y => l2c33_1, cin => l2c33_2, s => l3c33_3, cout => l3c34_0);
fulladder273: full_adder port map(x => l2c33_3, y => l2c33_4, cin => l2c33_5, s => l3c33_4, cout => l3c34_1);
fulladder274: full_adder port map(x => l2c33_6, y => l2c33_7, cin => l2c33_8, s => l3c33_5, cout => l3c34_2);
fulladder275: full_adder port map(x => l2c34_0, y => l2c34_1, cin => l2c34_2, s => l3c34_3, cout => l3c35_0);
fulladder276: full_adder port map(x => l2c34_3, y => l2c34_4, cin => l2c34_5, s => l3c34_4, cout => l3c35_1);
fulladder277: full_adder port map(x => l2c34_6, y => l2c34_7, cin => l2c34_8, s => l3c34_5, cout => l3c35_2);
fulladder278: full_adder port map(x => l2c35_0, y => l2c35_1, cin => l2c35_2, s => l3c35_3, cout => l3c36_0);
fulladder279: full_adder port map(x => l2c35_3, y => l2c35_4, cin => l2c35_5, s => l3c35_4, cout => l3c36_1);
fulladder280: full_adder port map(x => l2c36_0, y => l2c36_1, cin => l2c36_2, s => l3c36_3, cout => l3c37_0);
fulladder281: full_adder port map(x => l2c36_3, y => l2c36_4, cin => l2c36_5, s => l3c36_4, cout => l3c37_1);
fulladder282: full_adder port map(x => l2c37_0, y => l2c37_1, cin => l2c37_2, s => l3c37_3, cout => l3c38_0);
fulladder283: full_adder port map(x => l2c37_3, y => l2c37_4, cin => l2c37_5, s => l3c37_4, cout => l3c38_1);
fulladder284: full_adder port map(x => l2c38_0, y => l2c38_1, cin => l2c38_2, s => l3c38_3, cout => l3c39_0);
fulladder285: full_adder port map(x => l2c38_3, y => l2c38_4, cin => l2c38_5, s => l3c38_4, cout => l3c39_1);
fulladder286: full_adder port map(x => l2c39_0, y => l2c39_1, cin => l2c39_2, s => l3c39_2, cout => l3c40_0);
fulladder287: full_adder port map(x => l2c39_3, y => l2c39_4, cin => l2c39_5, s => l3c39_3, cout => l3c40_1);
fulladder288: full_adder port map(x => l2c40_0, y => l2c40_1, cin => l2c40_2, s => l3c40_2, cout => l3c41_0);
fulladder289: full_adder port map(x => l2c40_3, y => l2c40_4, cin => l1c40_6, s => l3c40_3, cout => l3c41_1);
fulladder290: full_adder port map(x => l2c41_0, y => l2c41_1, cin => l2c41_2, s => l3c41_2, cout => l3c42_0);
fulladder291: full_adder port map(x => l2c42_0, y => l2c42_1, cin => l2c42_2, s => l3c42_1, cout => l3c43_0);
fulladder292: full_adder port map(x => l2c43_0, y => l2c43_1, cin => l2c43_2, s => l3c43_1, cout => l3c44_0);
fulladder293: full_adder port map(x => l3c5_0, y => l3c5_1, cin => l2c5_3, s => l4c5_1, cout => l4c6_0);
fulladder294: full_adder port map(x => l3c6_0, y => l3c6_1, cin => l3c6_2, s => l4c6_1, cout => l4c7_0);
fulladder295: full_adder port map(x => l3c7_0, y => l3c7_1, cin => l3c7_2, s => l4c7_1, cout => l4c8_0);
fulladder296: full_adder port map(x => l3c8_0, y => l3c8_1, cin => l3c8_2, s => l4c8_1, cout => l4c9_0);
fulladder297: full_adder port map(x => l3c9_0, y => l3c9_1, cin => l3c9_2, s => l4c9_1, cout => l4c10_0);
fulladder298: full_adder port map(x => l3c10_0, y => l3c10_1, cin => l3c10_2, s => l4c10_2, cout => l4c11_0);
fulladder299: full_adder port map(x => l3c11_0, y => l3c11_1, cin => l3c11_2, s => l4c11_2, cout => l4c12_0);
fulladder300: full_adder port map(x => l3c12_0, y => l3c12_1, cin => l3c12_2, s => l4c12_2, cout => l4c13_0);
fulladder301: full_adder port map(x => l3c12_3, y => l3c12_4, cin => l3c12_5, s => l4c12_3, cout => l4c13_1);
fulladder302: full_adder port map(x => l3c13_0, y => l3c13_1, cin => l3c13_2, s => l4c13_2, cout => l4c14_0);
fulladder303: full_adder port map(x => l3c13_3, y => l3c13_4, cin => l3c13_5, s => l4c13_3, cout => l4c14_1);
fulladder304: full_adder port map(x => l3c14_0, y => l3c14_1, cin => l3c14_2, s => l4c14_2, cout => l4c15_0);
fulladder305: full_adder port map(x => l3c14_3, y => l3c14_4, cin => l3c14_5, s => l4c14_3, cout => l4c15_1);
fulladder306: full_adder port map(x => l3c15_0, y => l3c15_1, cin => l3c15_2, s => l4c15_2, cout => l4c16_0);
fulladder307: full_adder port map(x => l3c15_3, y => l3c15_4, cin => l3c15_5, s => l4c15_3, cout => l4c16_1);
fulladder308: full_adder port map(x => l3c16_0, y => l3c16_1, cin => l3c16_2, s => l4c16_2, cout => l4c17_0);
fulladder309: full_adder port map(x => l3c16_3, y => l3c16_4, cin => l3c16_5, s => l4c16_3, cout => l4c17_1);
fulladder310: full_adder port map(x => l3c17_0, y => l3c17_1, cin => l3c17_2, s => l4c17_3, cout => l4c18_0);
fulladder311: full_adder port map(x => l3c17_3, y => l3c17_4, cin => l3c17_5, s => l4c17_4, cout => l4c18_1);
fulladder312: full_adder port map(x => l3c18_0, y => l3c18_1, cin => l3c18_2, s => l4c18_3, cout => l4c19_0);
fulladder313: full_adder port map(x => l3c18_3, y => l3c18_4, cin => l3c18_5, s => l4c18_4, cout => l4c19_1);
fulladder314: full_adder port map(x => l3c18_6, y => l3c18_7, cin => l1c18_18, s => l4c18_5, cout => l4c19_2);
fulladder315: full_adder port map(x => l3c19_0, y => l3c19_1, cin => l3c19_2, s => l4c19_3, cout => l4c20_0);
fulladder316: full_adder port map(x => l3c19_3, y => l3c19_4, cin => l3c19_5, s => l4c19_4, cout => l4c20_1);
fulladder317: full_adder port map(x => l3c19_6, y => l3c19_7, cin => l2c19_12, s => l4c19_5, cout => l4c20_2);
fulladder318: full_adder port map(x => l3c20_0, y => l3c20_1, cin => l3c20_2, s => l4c20_3, cout => l4c21_0);
fulladder319: full_adder port map(x => l3c20_3, y => l3c20_4, cin => l3c20_5, s => l4c20_4, cout => l4c21_1);
fulladder320: full_adder port map(x => l3c20_6, y => l3c20_7, cin => l3c20_8, s => l4c20_5, cout => l4c21_2);
fulladder321: full_adder port map(x => l3c21_0, y => l3c21_1, cin => l3c21_2, s => l4c21_3, cout => l4c22_0);
fulladder322: full_adder port map(x => l3c21_3, y => l3c21_4, cin => l3c21_5, s => l4c21_4, cout => l4c22_1);
fulladder323: full_adder port map(x => l3c21_6, y => l3c21_7, cin => l3c21_8, s => l4c21_5, cout => l4c22_2);
fulladder324: full_adder port map(x => l3c22_0, y => l3c22_1, cin => l3c22_2, s => l4c22_3, cout => l4c23_0);
fulladder325: full_adder port map(x => l3c22_3, y => l3c22_4, cin => l3c22_5, s => l4c22_4, cout => l4c23_1);
fulladder326: full_adder port map(x => l3c22_6, y => l3c22_7, cin => l3c22_8, s => l4c22_5, cout => l4c23_2);
fulladder327: full_adder port map(x => l3c23_0, y => l3c23_1, cin => l3c23_2, s => l4c23_3, cout => l4c24_0);
fulladder328: full_adder port map(x => l3c23_3, y => l3c23_4, cin => l3c23_5, s => l4c23_4, cout => l4c24_1);
fulladder329: full_adder port map(x => l3c23_6, y => l3c23_7, cin => l3c23_8, s => l4c23_5, cout => l4c24_2);
fulladder330: full_adder port map(x => l3c24_0, y => l3c24_1, cin => l3c24_2, s => l4c24_4, cout => l4c25_0);
fulladder331: full_adder port map(x => l3c24_3, y => l3c24_4, cin => l3c24_5, s => l4c24_5, cout => l4c25_1);
fulladder332: full_adder port map(x => l3c24_6, y => l3c24_7, cin => l3c24_8, s => l4c24_6, cout => l4c25_2);
fulladder333: full_adder port map(x => l3c25_0, y => l3c25_1, cin => l3c25_2, s => l4c25_4, cout => l4c26_0);
fulladder334: full_adder port map(x => l3c25_3, y => l3c25_4, cin => l3c25_5, s => l4c25_5, cout => l4c26_1);
fulladder335: full_adder port map(x => l3c25_6, y => l3c25_7, cin => l3c25_8, s => l4c25_6, cout => l4c26_2);
fulladder336: full_adder port map(x => l3c26_0, y => l3c26_1, cin => l3c26_2, s => l4c26_4, cout => l4c27_0);
fulladder337: full_adder port map(x => l3c26_3, y => l3c26_4, cin => l3c26_5, s => l4c26_5, cout => l4c27_1);
fulladder338: full_adder port map(x => l3c26_6, y => l3c26_7, cin => l3c26_8, s => l4c26_6, cout => l4c27_2);
fulladder339: full_adder port map(x => l3c27_0, y => l3c27_1, cin => l3c27_2, s => l4c27_3, cout => l4c28_0);
fulladder340: full_adder port map(x => l3c27_3, y => l3c27_4, cin => l3c27_5, s => l4c27_4, cout => l4c28_1);
fulladder341: full_adder port map(x => l3c27_6, y => l3c27_7, cin => l3c27_8, s => l4c27_5, cout => l4c28_2);
fulladder342: full_adder port map(x => l3c28_0, y => l3c28_1, cin => l3c28_2, s => l4c28_3, cout => l4c29_0);
fulladder343: full_adder port map(x => l3c28_3, y => l3c28_4, cin => l3c28_5, s => l4c28_4, cout => l4c29_1);
fulladder344: full_adder port map(x => l3c28_6, y => l3c28_7, cin => l3c28_8, s => l4c28_5, cout => l4c29_2);
fulladder345: full_adder port map(x => l3c29_0, y => l3c29_1, cin => l3c29_2, s => l4c29_3, cout => l4c30_0);
fulladder346: full_adder port map(x => l3c29_3, y => l3c29_4, cin => l3c29_5, s => l4c29_4, cout => l4c30_1);
fulladder347: full_adder port map(x => l3c29_6, y => l3c29_7, cin => l3c29_8, s => l4c29_5, cout => l4c30_2);
fulladder348: full_adder port map(x => l3c30_0, y => l3c30_1, cin => l3c30_2, s => l4c30_3, cout => l4c31_0);
fulladder349: full_adder port map(x => l3c30_3, y => l3c30_4, cin => l3c30_5, s => l4c30_4, cout => l4c31_1);
fulladder350: full_adder port map(x => l3c31_0, y => l3c31_1, cin => l3c31_2, s => l4c31_3, cout => l4c32_0);
fulladder351: full_adder port map(x => l3c31_3, y => l3c31_4, cin => l3c31_5, s => l4c31_4, cout => l4c32_1);
fulladder352: full_adder port map(x => l3c32_0, y => l3c32_1, cin => l3c32_2, s => l4c32_3, cout => l4c33_0);
fulladder353: full_adder port map(x => l3c32_3, y => l3c32_4, cin => l3c32_5, s => l4c32_4, cout => l4c33_1);
fulladder354: full_adder port map(x => l3c33_0, y => l3c33_1, cin => l3c33_2, s => l4c33_3, cout => l4c34_0);
fulladder355: full_adder port map(x => l3c33_3, y => l3c33_4, cin => l3c33_5, s => l4c33_4, cout => l4c34_1);
fulladder356: full_adder port map(x => l3c34_0, y => l3c34_1, cin => l3c34_2, s => l4c34_2, cout => l4c35_0);
fulladder357: full_adder port map(x => l3c34_3, y => l3c34_4, cin => l3c34_5, s => l4c34_3, cout => l4c35_1);
fulladder358: full_adder port map(x => l3c35_0, y => l3c35_1, cin => l3c35_2, s => l4c35_2, cout => l4c36_0);
fulladder359: full_adder port map(x => l3c35_3, y => l3c35_4, cin => l3c35_5, s => l4c35_3, cout => l4c36_1);
fulladder360: full_adder port map(x => l3c36_0, y => l3c36_1, cin => l3c36_2, s => l4c36_2, cout => l4c37_0);
fulladder361: full_adder port map(x => l3c36_3, y => l3c36_4, cin => l3c36_5, s => l4c36_3, cout => l4c37_1);
fulladder362: full_adder port map(x => l3c37_0, y => l3c37_1, cin => l3c37_2, s => l4c37_2, cout => l4c38_0);
fulladder363: full_adder port map(x => l3c37_3, y => l3c37_4, cin => l3c37_5, s => l4c37_3, cout => l4c38_1);
fulladder364: full_adder port map(x => l3c38_0, y => l3c38_1, cin => l3c38_2, s => l4c38_2, cout => l4c39_0);
fulladder365: full_adder port map(x => l3c39_0, y => l3c39_1, cin => l3c39_2, s => l4c39_2, cout => l4c40_0);
fulladder366: full_adder port map(x => l3c40_0, y => l3c40_1, cin => l3c40_2, s => l4c40_1, cout => l4c41_0);
fulladder367: full_adder port map(x => l3c41_0, y => l3c41_1, cin => l3c41_2, s => l4c41_1, cout => l4c42_0);
fulladder368: full_adder port map(x => l3c42_0, y => l3c42_1, cin => l2c42_3, s => l4c42_1, cout => l4c43_0);
fulladder369: full_adder port map(x => l3c43_0, y => l3c43_1, cin => l1c43_3, s => l4c43_1, cout => l4c44_0);
fulladder370: full_adder port map(x => l4c7_0, y => l4c7_1, cin => l3c7_3, s => l5c7_1, cout => l5c8_0);
fulladder371: full_adder port map(x => l4c8_0, y => l4c8_1, cin => l3c8_3, s => l5c8_1, cout => l5c9_0);
fulladder372: full_adder port map(x => l4c9_0, y => l4c9_1, cin => l4c9_2, s => l5c9_1, cout => l5c10_0);
fulladder373: full_adder port map(x => l4c10_0, y => l4c10_1, cin => l4c10_2, s => l5c10_1, cout => l5c11_0);
fulladder374: full_adder port map(x => l4c11_0, y => l4c11_1, cin => l4c11_2, s => l5c11_1, cout => l5c12_0);
fulladder375: full_adder port map(x => l4c12_0, y => l4c12_1, cin => l4c12_2, s => l5c12_1, cout => l5c13_0);
fulladder376: full_adder port map(x => l4c13_0, y => l4c13_1, cin => l4c13_2, s => l5c13_1, cout => l5c14_0);
fulladder377: full_adder port map(x => l4c14_0, y => l4c14_1, cin => l4c14_2, s => l5c14_1, cout => l5c15_0);
fulladder378: full_adder port map(x => l4c15_0, y => l4c15_1, cin => l4c15_2, s => l5c15_2, cout => l5c16_0);
fulladder379: full_adder port map(x => l4c16_0, y => l4c16_1, cin => l4c16_2, s => l5c16_2, cout => l5c17_0);
fulladder380: full_adder port map(x => l4c17_0, y => l4c17_1, cin => l4c17_2, s => l5c17_2, cout => l5c18_0);
fulladder381: full_adder port map(x => l4c17_3, y => l4c17_4, cin => l4c17_5, s => l5c17_3, cout => l5c18_1);
fulladder382: full_adder port map(x => l4c18_0, y => l4c18_1, cin => l4c18_2, s => l5c18_2, cout => l5c19_0);
fulladder383: full_adder port map(x => l4c18_3, y => l4c18_4, cin => l4c18_5, s => l5c18_3, cout => l5c19_1);
fulladder384: full_adder port map(x => l4c19_0, y => l4c19_1, cin => l4c19_2, s => l5c19_2, cout => l5c20_0);
fulladder385: full_adder port map(x => l4c19_3, y => l4c19_4, cin => l4c19_5, s => l5c19_3, cout => l5c20_1);
fulladder386: full_adder port map(x => l4c20_0, y => l4c20_1, cin => l4c20_2, s => l5c20_2, cout => l5c21_0);
fulladder387: full_adder port map(x => l4c20_3, y => l4c20_4, cin => l4c20_5, s => l5c20_3, cout => l5c21_1);
fulladder388: full_adder port map(x => l4c21_0, y => l4c21_1, cin => l4c21_2, s => l5c21_2, cout => l5c22_0);
fulladder389: full_adder port map(x => l4c21_3, y => l4c21_4, cin => l4c21_5, s => l5c21_3, cout => l5c22_1);
fulladder390: full_adder port map(x => l4c22_0, y => l4c22_1, cin => l4c22_2, s => l5c22_2, cout => l5c23_0);
fulladder391: full_adder port map(x => l4c22_3, y => l4c22_4, cin => l4c22_5, s => l5c22_3, cout => l5c23_1);
fulladder392: full_adder port map(x => l4c23_0, y => l4c23_1, cin => l4c23_2, s => l5c23_2, cout => l5c24_0);
fulladder393: full_adder port map(x => l4c23_3, y => l4c23_4, cin => l4c23_5, s => l5c23_3, cout => l5c24_1);
fulladder394: full_adder port map(x => l4c24_0, y => l4c24_1, cin => l4c24_2, s => l5c24_2, cout => l5c25_0);
fulladder395: full_adder port map(x => l4c24_3, y => l4c24_4, cin => l4c24_5, s => l5c24_3, cout => l5c25_1);
fulladder396: full_adder port map(x => l4c25_0, y => l4c25_1, cin => l4c25_2, s => l5c25_3, cout => l5c26_0);
fulladder397: full_adder port map(x => l4c25_3, y => l4c25_4, cin => l4c25_5, s => l5c25_4, cout => l5c26_1);
fulladder398: full_adder port map(x => l4c26_0, y => l4c26_1, cin => l4c26_2, s => l5c26_3, cout => l5c27_0);
fulladder399: full_adder port map(x => l4c26_3, y => l4c26_4, cin => l4c26_5, s => l5c26_4, cout => l5c27_1);
fulladder400: full_adder port map(x => l4c27_0, y => l4c27_1, cin => l4c27_2, s => l5c27_3, cout => l5c28_0);
fulladder401: full_adder port map(x => l4c27_3, y => l4c27_4, cin => l4c27_5, s => l5c27_4, cout => l5c28_1);
fulladder402: full_adder port map(x => l4c28_0, y => l4c28_1, cin => l4c28_2, s => l5c28_2, cout => l5c29_0);
fulladder403: full_adder port map(x => l4c28_3, y => l4c28_4, cin => l4c28_5, s => l5c28_3, cout => l5c29_1);
fulladder404: full_adder port map(x => l4c29_0, y => l4c29_1, cin => l4c29_2, s => l5c29_2, cout => l5c30_0);
fulladder405: full_adder port map(x => l4c29_3, y => l4c29_4, cin => l4c29_5, s => l5c29_3, cout => l5c30_1);
fulladder406: full_adder port map(x => l4c30_0, y => l4c30_1, cin => l4c30_2, s => l5c30_2, cout => l5c31_0);
fulladder407: full_adder port map(x => l4c30_3, y => l4c30_4, cin => l4c30_5, s => l5c30_3, cout => l5c31_1);
fulladder408: full_adder port map(x => l4c31_0, y => l4c31_1, cin => l4c31_2, s => l5c31_2, cout => l5c32_0);
fulladder409: full_adder port map(x => l4c31_3, y => l4c31_4, cin => l4c31_5, s => l5c31_3, cout => l5c32_1);
fulladder410: full_adder port map(x => l4c32_0, y => l4c32_1, cin => l4c32_2, s => l5c32_2, cout => l5c33_0);
fulladder411: full_adder port map(x => l4c32_3, y => l4c32_4, cin => l4c32_5, s => l5c32_3, cout => l5c33_1);
fulladder412: full_adder port map(x => l4c33_0, y => l4c33_1, cin => l4c33_2, s => l5c33_2, cout => l5c34_0);
fulladder413: full_adder port map(x => l4c33_3, y => l4c33_4, cin => l2c33_9, s => l5c33_3, cout => l5c34_1);
fulladder414: full_adder port map(x => l4c34_0, y => l4c34_1, cin => l4c34_2, s => l5c34_2, cout => l5c35_0);
fulladder415: full_adder port map(x => l4c35_0, y => l4c35_1, cin => l4c35_2, s => l5c35_2, cout => l5c36_0);
fulladder416: full_adder port map(x => l4c36_0, y => l4c36_1, cin => l4c36_2, s => l5c36_1, cout => l5c37_0);
fulladder417: full_adder port map(x => l4c37_0, y => l4c37_1, cin => l4c37_2, s => l5c37_1, cout => l5c38_0);
fulladder418: full_adder port map(x => l4c38_0, y => l4c38_1, cin => l4c38_2, s => l5c38_1, cout => l5c39_0);
fulladder419: full_adder port map(x => l4c39_0, y => l4c39_1, cin => l4c39_2, s => l5c39_1, cout => l5c40_0);
fulladder420: full_adder port map(x => l4c40_0, y => l4c40_1, cin => l3c40_3, s => l5c40_1, cout => l5c41_0);
fulladder421: full_adder port map(x => l4c41_0, y => l4c41_1, cin => l2c41_3, s => l5c41_1, cout => l5c42_0);
fulladder422: full_adder port map(x => l5c10_0, y => l5c10_1, cin => l4c10_3, s => l6c10_1, cout => l6c11_0);
fulladder423: full_adder port map(x => l5c11_0, y => l5c11_1, cin => l4c11_3, s => l6c11_1, cout => l6c12_0);
fulladder424: full_adder port map(x => l5c12_0, y => l5c12_1, cin => l4c12_3, s => l6c12_1, cout => l6c13_0);
fulladder425: full_adder port map(x => l5c13_0, y => l5c13_1, cin => l4c13_3, s => l6c13_1, cout => l6c14_0);
fulladder426: full_adder port map(x => l5c14_0, y => l5c14_1, cin => l5c14_2, s => l6c14_1, cout => l6c15_0);
fulladder427: full_adder port map(x => l5c15_0, y => l5c15_1, cin => l5c15_2, s => l6c15_1, cout => l6c16_0);
fulladder428: full_adder port map(x => l5c16_0, y => l5c16_1, cin => l5c16_2, s => l6c16_1, cout => l6c17_0);
fulladder429: full_adder port map(x => l5c17_0, y => l5c17_1, cin => l5c17_2, s => l6c17_1, cout => l6c18_0);
fulladder430: full_adder port map(x => l5c18_0, y => l5c18_1, cin => l5c18_2, s => l6c18_1, cout => l6c19_0);
fulladder431: full_adder port map(x => l5c19_0, y => l5c19_1, cin => l5c19_2, s => l6c19_1, cout => l6c20_0);
fulladder432: full_adder port map(x => l5c20_0, y => l5c20_1, cin => l5c20_2, s => l6c20_1, cout => l6c21_0);
fulladder433: full_adder port map(x => l5c21_0, y => l5c21_1, cin => l5c21_2, s => l6c21_1, cout => l6c22_0);
fulladder434: full_adder port map(x => l5c22_0, y => l5c22_1, cin => l5c22_2, s => l6c22_2, cout => l6c23_0);
fulladder435: full_adder port map(x => l5c23_0, y => l5c23_1, cin => l5c23_2, s => l6c23_2, cout => l6c24_0);
fulladder436: full_adder port map(x => l5c24_0, y => l5c24_1, cin => l5c24_2, s => l6c24_2, cout => l6c25_0);
fulladder437: full_adder port map(x => l5c25_0, y => l5c25_1, cin => l5c25_2, s => l6c25_2, cout => l6c26_0);
fulladder438: full_adder port map(x => l5c25_3, y => l5c25_4, cin => l5c25_5, s => l6c25_3, cout => l6c26_1);
fulladder439: full_adder port map(x => l5c26_0, y => l5c26_1, cin => l5c26_2, s => l6c26_2, cout => l6c27_0);
fulladder440: full_adder port map(x => l5c26_3, y => l5c26_4, cin => l5c26_5, s => l6c26_3, cout => l6c27_1);
fulladder441: full_adder port map(x => l5c27_0, y => l5c27_1, cin => l5c27_2, s => l6c27_2, cout => l6c28_0);
fulladder442: full_adder port map(x => l5c27_3, y => l5c27_4, cin => l3c27_9, s => l6c27_3, cout => l6c28_1);
fulladder443: full_adder port map(x => l5c28_0, y => l5c28_1, cin => l5c28_2, s => l6c28_2, cout => l6c29_0);
fulladder444: full_adder port map(x => l5c29_0, y => l5c29_1, cin => l5c29_2, s => l6c29_2, cout => l6c30_0);
fulladder445: full_adder port map(x => l5c30_0, y => l5c30_1, cin => l5c30_2, s => l6c30_1, cout => l6c31_0);
fulladder446: full_adder port map(x => l5c31_0, y => l5c31_1, cin => l5c31_2, s => l6c31_1, cout => l6c32_0);
fulladder447: full_adder port map(x => l5c32_0, y => l5c32_1, cin => l5c32_2, s => l6c32_1, cout => l6c33_0);
fulladder448: full_adder port map(x => l5c33_0, y => l5c33_1, cin => l5c33_2, s => l6c33_1, cout => l6c34_0);
fulladder449: full_adder port map(x => l5c34_0, y => l5c34_1, cin => l5c34_2, s => l6c34_1, cout => l6c35_0);
fulladder450: full_adder port map(x => l5c35_0, y => l5c35_1, cin => l5c35_2, s => l6c35_1, cout => l6c36_0);
fulladder451: full_adder port map(x => l5c36_0, y => l5c36_1, cin => l4c36_3, s => l6c36_1, cout => l6c37_0);
fulladder452: full_adder port map(x => l5c37_0, y => l5c37_1, cin => l4c37_3, s => l6c37_1, cout => l6c38_0);
fulladder453: full_adder port map(x => l5c38_0, y => l5c38_1, cin => l4c38_3, s => l6c38_1, cout => l6c39_0);
fulladder454: full_adder port map(x => l5c39_0, y => l5c39_1, cin => l3c39_3, s => l6c39_1, cout => l6c40_0);
fulladder455: full_adder port map(x => l6c15_0, y => l6c15_1, cin => l5c15_3, s => l7c15_1, cout => l7c16_0);
fulladder456: full_adder port map(x => l6c16_0, y => l6c16_1, cin => l5c16_3, s => l7c16_1, cout => l7c17_0);
fulladder457: full_adder port map(x => l6c17_0, y => l6c17_1, cin => l5c17_3, s => l7c17_1, cout => l7c18_0);
fulladder458: full_adder port map(x => l6c18_0, y => l6c18_1, cin => l5c18_3, s => l7c18_1, cout => l7c19_0);
fulladder459: full_adder port map(x => l6c19_0, y => l6c19_1, cin => l5c19_3, s => l7c19_1, cout => l7c20_0);
fulladder460: full_adder port map(x => l6c20_0, y => l6c20_1, cin => l5c20_3, s => l7c20_1, cout => l7c21_0);
fulladder461: full_adder port map(x => l6c21_0, y => l6c21_1, cin => l6c21_2, s => l7c21_1, cout => l7c22_0);
fulladder462: full_adder port map(x => l6c22_0, y => l6c22_1, cin => l6c22_2, s => l7c22_1, cout => l7c23_0);
fulladder463: full_adder port map(x => l6c23_0, y => l6c23_1, cin => l6c23_2, s => l7c23_1, cout => l7c24_0);
fulladder464: full_adder port map(x => l6c24_0, y => l6c24_1, cin => l6c24_2, s => l7c24_1, cout => l7c25_0);
fulladder465: full_adder port map(x => l6c25_0, y => l6c25_1, cin => l6c25_2, s => l7c25_1, cout => l7c26_0);
fulladder466: full_adder port map(x => l6c26_0, y => l6c26_1, cin => l6c26_2, s => l7c26_1, cout => l7c27_0);
fulladder467: full_adder port map(x => l6c27_0, y => l6c27_1, cin => l6c27_2, s => l7c27_1, cout => l7c28_0);
fulladder468: full_adder port map(x => l6c28_0, y => l6c28_1, cin => l6c28_2, s => l7c28_1, cout => l7c29_0);
fulladder469: full_adder port map(x => l6c29_0, y => l6c29_1, cin => l6c29_2, s => l7c29_1, cout => l7c30_0);
fulladder470: full_adder port map(x => l6c30_0, y => l6c30_1, cin => l5c30_3, s => l7c30_1, cout => l7c31_0);
fulladder471: full_adder port map(x => l6c31_0, y => l6c31_1, cin => l5c31_3, s => l7c31_1, cout => l7c32_0);
fulladder472: full_adder port map(x => l6c32_0, y => l6c32_1, cin => l5c32_3, s => l7c32_1, cout => l7c33_0);
fulladder473: full_adder port map(x => l6c33_0, y => l6c33_1, cin => l5c33_3, s => l7c33_1, cout => l7c34_0);
fulladder474: full_adder port map(x => l6c34_0, y => l6c34_1, cin => l5c34_3, s => l7c34_1, cout => l7c35_0);
fulladder475: full_adder port map(x => l6c35_0, y => l6c35_1, cin => l4c35_3, s => l7c35_1, cout => l7c36_0);
fulladder476: full_adder port map(x => l7c22_0, y => l7c22_1, cin => l6c22_3, s => l8c22_1, cout => l8c23_0);
fulladder477: full_adder port map(x => l7c23_0, y => l7c23_1, cin => l6c23_3, s => l8c23_1, cout => l8c24_0);
fulladder478: full_adder port map(x => l7c24_0, y => l7c24_1, cin => l6c24_3, s => l8c24_1, cout => l8c25_0);
fulladder479: full_adder port map(x => l7c25_0, y => l7c25_1, cin => l6c25_3, s => l8c25_1, cout => l8c26_0);
fulladder480: full_adder port map(x => l7c26_0, y => l7c26_1, cin => l6c26_3, s => l8c26_1, cout => l8c27_0);
fulladder481: full_adder port map(x => l7c27_0, y => l7c27_1, cin => l6c27_3, s => l8c27_1, cout => l8c28_0);
fulladder482: full_adder port map(x => l7c28_0, y => l7c28_1, cin => l6c28_3, s => l8c28_1, cout => l8c29_0);
fulladder483: full_adder port map(x => l7c29_0, y => l7c29_1, cin => l5c29_3, s => l8c29_1, cout => l8c30_0);

final_x <= l8c47_0 & l8c46_0 & l8c45_0 & l8c44_0 & l8c43_0 & l8c42_0 & l8c41_0 & l8c40_0 & l8c39_0 & l8c38_0 & l8c37_0 & l8c36_0 & l8c35_0 & l8c34_0 & l8c33_0 & l8c32_0 & l8c31_0 & l8c30_0 & l8c29_0 & l8c28_0 & l8c27_0 & l8c26_0 & l8c25_0 & l8c24_0 & l8c23_0 & l8c22_0 & l8c21_0 & l8c20_0 & l8c19_0 & l8c18_0 & l8c17_0 & l8c16_0 & l8c15_0 & l8c14_0 & l8c13_0 & l8c12_0 & l8c11_0 & l8c10_0 & l8c9_0 & l8c8_0 & l8c7_0 & l7c6_0 & l6c5_0 & l5c4_0 & l4c3_0 & l3c2_0 & l2c1_0 & l1c0_0;
final_y <= l8c47_1 & l8c46_1 & l8c45_1 & l8c44_1 & l8c43_1 & l8c42_1 & l8c41_1 & l8c40_1 & l8c39_1 & l8c38_1 & l8c37_1 & l8c36_1 & l8c35_1 & l8c34_1 & l8c33_1 & l8c32_1 & l8c31_1 & l8c30_1 & l8c29_1 & l8c28_1 & l8c27_1 & l8c26_1 & l8c25_1 & l8c24_1 & l8c23_1 & l8c22_1 & l8c21_1 & l8c20_1 & l8c19_1 & l8c18_1 & l8c17_1 & l8c16_1 & l8c15_1 & l8c14_1 & l8c13_1 & l8c12_1 & l8c11_1 & l8c10_1 & l8c9_1 & l8c8_1 & b"0" & b"0" & b"0" & b"0" & b"0" & b"0" & b"0" & b"0";
final_adder: carry_lookahead_adder_48 port map(final_x, final_y, '0', p);

end arch;